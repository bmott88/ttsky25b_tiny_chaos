magic
tech sky130A
timestamp 1762404587
<< nwell >>
rect 2539 535 2670 1847
rect 2539 -3167 2670 -543
rect 2351 -5225 2670 -4245
rect 1069 -5557 2688 -5225
<< pwell >>
rect -1535 1524 -22 1847
rect -380 -3541 -22 1524
rect 2539 -543 2670 535
rect 41 -3541 2826 -3167
rect -380 -4245 2826 -3541
rect 5231 -3207 5789 1847
rect -380 -4272 1173 -4245
rect -380 -5195 1168 -4272
rect -1535 -5196 1168 -5195
rect -1535 -5557 1069 -5196
rect 5231 -5557 7685 -3207
rect 5469 -5558 5789 -5557
<< metal1 >>
rect -22 1913 7685 1950
rect -22 1876 2791 1913
rect 2977 1912 7685 1913
rect 2977 1876 4764 1912
rect -22 1859 4764 1876
rect 5149 1859 7685 1912
rect -22 1821 7685 1859
rect -22 1809 4998 1821
rect -1535 1638 -380 1695
rect -1535 1533 -1456 1638
rect -479 1533 -380 1638
rect -22 1550 302 1809
rect 2215 1733 2995 1809
rect 2215 1696 2767 1733
rect 2953 1696 2995 1733
rect 2215 1550 2995 1696
rect 4907 1735 4998 1809
rect 5137 1807 7685 1821
rect 5137 1735 5231 1807
rect 4907 1550 5231 1735
rect -1535 1479 -380 1533
rect 2371 1488 2444 1500
rect -679 705 -463 1441
rect -284 1323 -211 1335
rect -284 1144 -272 1323
rect -226 1252 -211 1323
rect 2371 1309 2383 1488
rect 2429 1333 2444 1488
rect 5192 1448 5266 1468
rect 5701 1459 5813 1476
rect 5701 1448 5724 1459
rect 5192 1447 5724 1448
rect 5192 1407 5209 1447
rect 5244 1408 5724 1447
rect 5244 1407 5266 1408
rect 5192 1387 5266 1407
rect 5701 1399 5724 1408
rect 5786 1399 5813 1459
rect 7634 1408 7680 1448
rect 5701 1379 5813 1399
rect 2429 1309 2712 1333
rect 2371 1297 2712 1309
rect 2670 1252 2712 1297
rect -226 1226 146 1252
rect 2670 1226 2838 1252
rect -226 1144 -211 1226
rect -284 1132 -211 1144
rect 5585 809 5808 828
rect 5585 761 5603 809
rect 5641 788 5808 809
rect 7634 788 7680 828
rect 5641 761 5659 788
rect -679 594 -610 705
rect -532 594 -463 705
rect 2568 751 2632 759
rect -1452 -53 -1236 69
rect -1452 -330 -1391 -53
rect -1313 -330 -1236 -53
rect -1452 -1190 -1236 -330
rect -679 -504 -463 594
rect -267 631 1282 657
rect -267 -93 -205 631
rect 2568 529 2578 751
rect 2621 657 2632 751
rect 5585 741 5659 761
rect 2621 631 3974 657
rect 2621 529 2632 631
rect 2568 521 2632 529
rect -22 94 570 274
rect -328 -129 -146 -93
rect -328 -264 -305 -129
rect -178 -264 -146 -129
rect -328 -294 -146 -264
rect -22 -103 98 94
rect 397 34 570 94
rect 1947 91 3262 274
rect 1947 34 2046 91
rect 397 -42 2046 34
rect 397 -103 570 -42
rect -22 -282 570 -103
rect 1947 -83 2046 -42
rect 2221 34 3262 91
rect 4639 34 5231 274
rect 2221 -42 5231 34
rect 2221 -83 3262 -42
rect 1947 -282 3262 -83
rect 4639 -282 5231 -42
rect 5606 1 5812 14
rect 5606 -52 5611 1
rect 5796 -52 5812 1
rect 7634 -50 7680 -10
rect 5606 -63 5812 -52
rect 5606 -64 5765 -63
rect 2571 -550 2635 -542
rect -679 -639 -463 -617
rect -679 -665 1282 -639
rect -1452 -1421 -1236 -1303
rect -1452 -1614 -1398 -1421
rect -1306 -1614 -1236 -1421
rect -1452 -2562 -1236 -1614
rect -679 -1876 -463 -665
rect 2571 -772 2581 -550
rect 2624 -639 2635 -550
rect 5512 -609 5623 -598
rect 5192 -625 5269 -614
rect 2624 -665 3974 -639
rect 2624 -772 2635 -665
rect 5192 -672 5204 -625
rect 5254 -630 5269 -625
rect 5512 -630 5523 -609
rect 5254 -670 5523 -630
rect 5254 -672 5269 -670
rect 5192 -683 5269 -672
rect 5512 -690 5523 -670
rect 5609 -630 5623 -609
rect 5609 -670 5842 -630
rect 5609 -690 5623 -670
rect 5512 -700 5623 -690
rect 2571 -780 2635 -772
rect -280 -1171 -207 -1159
rect -280 -1350 -268 -1171
rect -222 -1234 -207 -1171
rect -222 -1260 146 -1234
rect 2665 -1260 2838 -1234
rect -222 -1350 -207 -1260
rect 2665 -1307 2689 -1260
rect -280 -1362 -207 -1350
rect 2379 -1319 2689 -1307
rect 2379 -1498 2391 -1319
rect 2437 -1325 2689 -1319
rect 2437 -1498 2452 -1325
rect 2379 -1510 2452 -1498
rect 5428 -1455 5614 -1437
rect 5428 -1511 5446 -1455
rect 5571 -1468 5614 -1455
rect 5571 -1508 5808 -1468
rect 5571 -1511 5614 -1508
rect 5428 -1532 5614 -1511
rect -22 -1817 302 -1558
rect 2214 -1698 2994 -1558
rect 2214 -1739 2754 -1698
rect 2933 -1739 2994 -1698
rect 2214 -1817 2994 -1739
rect 4907 -1756 5231 -1558
rect 4907 -1817 4972 -1756
rect -22 -1893 4972 -1817
rect -1452 -2983 -1236 -2675
rect -1452 -3173 -1373 -2983
rect -1301 -3173 -1236 -2983
rect -1452 -3934 -1236 -3173
rect -679 -3045 -463 -1989
rect -22 -2152 302 -1893
rect 2214 -1973 2994 -1893
rect 2214 -2014 2757 -1973
rect 2936 -2014 2994 -1973
rect 2214 -2152 2994 -2014
rect 4907 -1940 4972 -1893
rect 5156 -1940 5231 -1756
rect 4907 -2152 5231 -1940
rect 5549 -2085 5624 -2071
rect 5549 -2136 5563 -2085
rect 5611 -2088 5624 -2085
rect 5611 -2127 5802 -2088
rect 5611 -2128 5799 -2127
rect 5611 -2136 5624 -2128
rect 5549 -2153 5624 -2136
rect 2372 -2219 2445 -2207
rect -283 -2385 -210 -2373
rect -283 -2564 -271 -2385
rect -225 -2450 -210 -2385
rect 2372 -2398 2384 -2219
rect 2430 -2381 2445 -2219
rect 5567 -2234 5597 -2153
rect 5192 -2246 5597 -2234
rect 5192 -2300 5204 -2246
rect 5259 -2258 5597 -2246
rect 5259 -2300 5275 -2258
rect 5192 -2314 5275 -2300
rect 2430 -2398 2700 -2381
rect 2372 -2410 2700 -2398
rect 2666 -2450 2700 -2410
rect -225 -2476 146 -2450
rect 2666 -2476 2838 -2450
rect -225 -2564 -210 -2476
rect -283 -2576 -210 -2564
rect 5649 -2940 5799 -2926
rect 2569 -2952 2633 -2944
rect -679 -3071 1282 -3045
rect -679 -3248 -463 -3071
rect 2569 -3174 2579 -2952
rect 2622 -3045 2633 -2952
rect 5649 -3000 5662 -2940
rect 5727 -2966 5799 -2940
rect 5727 -3000 5745 -2966
rect 5649 -3014 5745 -3000
rect 2622 -3071 3974 -3045
rect 2622 -3174 2633 -3071
rect 2569 -3182 2633 -3174
rect 5789 -3279 7685 -3216
rect 6179 -3315 7332 -3279
rect 7573 -3315 7685 -3279
rect -679 -4268 -463 -3361
rect 6179 -3427 7685 -3315
rect 5789 -3428 7685 -3427
rect -22 -3613 570 -3428
rect -22 -3810 67 -3613
rect 366 -3668 570 -3613
rect 1947 -3593 3262 -3428
rect 1947 -3668 2035 -3593
rect 366 -3767 2035 -3668
rect 2210 -3668 3262 -3593
rect 4639 -3560 7685 -3428
rect 4639 -3668 5231 -3560
rect 2210 -3744 5231 -3668
rect 2210 -3767 3262 -3744
rect 366 -3810 3262 -3767
rect -22 -3878 3262 -3810
rect 2670 -3984 3262 -3878
rect 4639 -3984 5231 -3744
rect -679 -4414 -645 -4268
rect -532 -4414 -463 -4268
rect -679 -5306 -463 -4414
rect 2548 -4243 2621 -4232
rect 2548 -4464 2560 -4243
rect 2606 -4341 2621 -4243
rect 2606 -4367 3974 -4341
rect 2606 -4464 2621 -4367
rect 2548 -4476 2621 -4464
rect -287 -4834 -156 -4816
rect -287 -5031 -268 -4834
rect -185 -5031 -156 -4834
rect 2369 -4932 2577 -4915
rect 2369 -4970 2386 -4932
rect 2557 -4936 2577 -4932
rect 2557 -4962 2838 -4936
rect 2557 -4970 2577 -4962
rect 2369 -4983 2577 -4970
rect -287 -5049 -156 -5031
rect 688 -5191 890 -5159
rect 688 -5309 724 -5191
rect 853 -5294 890 -5191
rect 853 -5309 1201 -5294
rect -1535 -5389 -380 -5344
rect 688 -5380 1201 -5309
rect 2233 -5308 2337 -5293
rect 2233 -5373 2249 -5308
rect 2318 -5373 2337 -5308
rect 2233 -5386 2337 -5373
rect 2670 -5406 2994 -5260
rect 2670 -5442 2753 -5406
rect 2937 -5442 2994 -5406
rect 2670 -5454 2994 -5442
rect -22 -5519 2994 -5454
rect 4906 -5304 7683 -5260
rect 4906 -5306 6873 -5304
rect 4906 -5438 5979 -5306
rect 4906 -5519 4981 -5438
rect -22 -5555 4981 -5519
rect 5159 -5555 5979 -5438
rect -22 -5558 5979 -5555
rect 6123 -5558 6873 -5306
rect -22 -5560 6873 -5558
rect -22 -5596 2796 -5560
rect 2980 -5585 6873 -5560
rect 7061 -5585 7683 -5304
rect 2980 -5596 7683 -5585
rect -22 -5620 7683 -5596
rect -22 -5621 5231 -5620
<< via1 >>
rect 2791 1876 2977 1913
rect 4764 1859 5149 1912
rect -1456 1533 -479 1638
rect 2767 1696 2953 1733
rect 4998 1735 5137 1821
rect -272 1144 -226 1323
rect 2383 1309 2429 1488
rect 5209 1407 5244 1447
rect 5724 1399 5786 1459
rect 5603 761 5641 809
rect -610 594 -532 705
rect -1391 -330 -1313 -53
rect 2578 529 2621 751
rect -305 -264 -178 -129
rect 98 -103 397 94
rect 2046 -83 2221 91
rect 5611 -52 5796 1
rect -1398 -1614 -1306 -1421
rect 2581 -772 2624 -550
rect 5204 -672 5254 -625
rect 5523 -690 5609 -609
rect -268 -1350 -222 -1171
rect 2391 -1498 2437 -1319
rect 5446 -1511 5571 -1455
rect 2754 -1739 2933 -1698
rect -1373 -3173 -1301 -2983
rect 2757 -2014 2936 -1973
rect 4972 -1940 5156 -1756
rect 5563 -2136 5611 -2085
rect -271 -2564 -225 -2385
rect 2384 -2398 2430 -2219
rect 5204 -2300 5259 -2246
rect 2579 -3174 2622 -2952
rect 5662 -3000 5727 -2940
rect 7332 -3315 7573 -3279
rect 67 -3810 366 -3613
rect 2035 -3767 2210 -3593
rect -645 -4414 -532 -4268
rect 2560 -4464 2606 -4243
rect -268 -5031 -185 -4834
rect 2386 -4970 2557 -4932
rect 724 -5309 853 -5191
rect 2249 -5373 2318 -5308
rect 2753 -5442 2937 -5406
rect 4981 -5555 5159 -5438
rect 5979 -5558 6123 -5306
rect 2796 -5596 2980 -5560
rect 6873 -5585 7061 -5304
<< metal2 >>
rect 2774 1913 2997 1928
rect 686 1860 846 1878
rect 686 1804 703 1860
rect -22 1796 703 1804
rect 826 1804 846 1860
rect 2774 1876 2791 1913
rect 2977 1876 2997 1913
rect 2774 1859 2997 1876
rect 4743 1912 5182 1926
rect 4743 1859 4764 1912
rect 5149 1859 5182 1912
rect 4743 1840 5182 1859
rect 4961 1821 5182 1840
rect 826 1796 3963 1804
rect -22 1778 3963 1796
rect 2756 1733 2964 1741
rect 2756 1696 2767 1733
rect 2953 1696 2964 1733
rect 4961 1735 4998 1821
rect 5137 1735 5182 1821
rect 4961 1704 5182 1735
rect 2756 1689 2964 1696
rect -1483 1638 -447 1662
rect -1483 1533 -1456 1638
rect -479 1533 -447 1638
rect -1483 1509 -447 1533
rect 2371 1488 2444 1500
rect -284 1323 -211 1335
rect -284 1144 -272 1323
rect -226 1144 -211 1323
rect 2371 1309 2383 1488
rect 2429 1309 2444 1488
rect 2371 1297 2444 1309
rect -284 1132 -211 1144
rect -633 705 -513 720
rect -633 594 -610 705
rect -532 594 -513 705
rect -633 578 -513 594
rect 57 94 443 133
rect -1413 -53 -1289 -24
rect -1413 -330 -1391 -53
rect -1313 -163 -1289 -53
rect -328 -129 -146 -93
rect -328 -163 -305 -129
rect -1313 -227 -305 -163
rect -1313 -330 -1289 -227
rect -328 -264 -305 -227
rect -178 -264 -146 -129
rect 57 -103 98 94
rect 397 -103 443 94
rect 57 -132 443 -103
rect 2008 91 2260 127
rect 2008 -83 2046 91
rect 2221 -83 2260 91
rect 2500 54 2526 1648
rect 5192 1468 5218 1648
rect 5192 1447 5266 1468
rect 5192 1407 5209 1447
rect 5244 1407 5266 1447
rect 5192 1387 5266 1407
rect 5701 1459 5813 1476
rect 5701 1399 5724 1459
rect 5786 1399 5813 1459
rect 2568 751 2632 759
rect 2568 529 2578 751
rect 2621 529 2632 751
rect 2568 521 2632 529
rect 5192 196 5218 1387
rect 5701 1379 5813 1399
rect 5585 814 5750 828
rect 5585 809 5653 814
rect 5585 783 5603 809
rect 5521 761 5603 783
rect 5641 761 5653 809
rect 5521 753 5653 761
rect 5720 753 5750 814
rect 5521 741 5750 753
rect 5521 54 5562 741
rect 2500 20 5562 54
rect 2500 19 5521 20
rect 5576 1 5812 14
rect 5576 -28 5611 1
rect 2008 -114 2260 -83
rect 2500 -52 5611 -28
rect 5796 -52 5812 1
rect 2500 -63 5812 -52
rect -328 -294 -146 -264
rect -1413 -368 -1289 -330
rect -280 -1171 -207 -1159
rect -280 -1350 -268 -1171
rect -222 -1350 -207 -1171
rect -280 -1362 -207 -1350
rect 2379 -1319 2452 -1307
rect -1426 -1421 -1273 -1388
rect -1426 -1614 -1398 -1421
rect -1306 -1614 -1273 -1421
rect 2379 -1498 2391 -1319
rect 2437 -1498 2452 -1319
rect 2379 -1510 2452 -1498
rect -1426 -1638 -1273 -1614
rect 2500 -1656 2526 -63
rect 5576 -64 5736 -63
rect 2571 -550 2635 -542
rect 2571 -772 2581 -550
rect 2624 -772 2635 -550
rect 2571 -780 2635 -772
rect 5192 -614 5218 -204
rect 5512 -609 5623 -598
rect 5192 -625 5269 -614
rect 5192 -672 5204 -625
rect 5254 -672 5269 -625
rect 5192 -683 5269 -672
rect 5192 -1309 5218 -683
rect 5512 -690 5523 -609
rect 5609 -690 5623 -609
rect 5512 -700 5623 -690
rect 5428 -1455 5614 -1437
rect 5428 -1511 5446 -1455
rect 5584 -1511 5614 -1455
rect 5428 -1532 5614 -1511
rect 5192 -1656 5218 -1557
rect 2744 -1698 2946 -1689
rect 2744 -1739 2754 -1698
rect 2933 -1739 2946 -1698
rect 2744 -1752 2946 -1739
rect 4954 -1756 5186 -1725
rect -22 -1800 3963 -1786
rect -22 -1908 709 -1800
rect 824 -1908 3963 -1800
rect -22 -1923 3963 -1908
rect 4954 -1940 4972 -1756
rect 5156 -1940 5186 -1756
rect 2738 -1973 2953 -1963
rect 4954 -1970 5186 -1940
rect 2738 -2014 2757 -1973
rect 2936 -2014 2953 -1973
rect 2738 -2025 2953 -2014
rect 2372 -2219 2445 -2207
rect -283 -2385 -210 -2373
rect -283 -2564 -271 -2385
rect -225 -2564 -210 -2385
rect 2372 -2398 2384 -2219
rect 2430 -2398 2445 -2219
rect 2372 -2410 2445 -2398
rect -283 -2576 -210 -2564
rect -1402 -2983 -1274 -2966
rect -1402 -3173 -1373 -2983
rect -1301 -3173 -1274 -2983
rect -1402 -3200 -1274 -3173
rect 28 -3613 414 -3584
rect 28 -3810 67 -3613
rect 366 -3810 414 -3613
rect 2012 -3593 2239 -3563
rect 2012 -3767 2035 -3593
rect 2210 -3767 2239 -3593
rect 2500 -3684 2526 -2054
rect 5192 -2234 5218 -2054
rect 5192 -2246 5275 -2234
rect 5192 -2300 5204 -2246
rect 5259 -2300 5275 -2246
rect 5192 -2314 5275 -2300
rect 2569 -2952 2633 -2944
rect 2569 -3174 2579 -2952
rect 2622 -3174 2633 -2952
rect 2569 -3182 2633 -3174
rect 5192 -3506 5218 -2314
rect 5429 -3684 5472 -1532
rect 5549 -2085 5624 -2071
rect 5549 -2136 5563 -2085
rect 5611 -2136 5624 -2085
rect 5549 -2153 5624 -2136
rect 2500 -3720 5472 -3684
rect 5649 -2938 5745 -2927
rect 5649 -3001 5662 -2938
rect 5729 -3001 5745 -2938
rect 5649 -3014 5745 -3001
rect 2012 -3796 2239 -3767
rect 28 -3849 414 -3810
rect 5649 -3906 5693 -3014
rect 7323 -3277 7588 -3232
rect 7323 -3315 7332 -3277
rect 7573 -3315 7588 -3277
rect 7323 -3329 7588 -3315
rect 5190 -3932 5693 -3906
rect -664 -4268 -503 -4242
rect -664 -4414 -645 -4268
rect -532 -4301 -503 -4268
rect 2548 -4243 2621 -4232
rect 2548 -4301 2560 -4243
rect -532 -4372 2560 -4301
rect -532 -4414 -503 -4372
rect -664 -4436 -503 -4414
rect 2548 -4464 2560 -4372
rect 2606 -4464 2621 -4243
rect 2548 -4476 2621 -4464
rect -287 -4834 -156 -4816
rect -287 -5031 -268 -4834
rect -185 -4915 -156 -4834
rect -185 -4932 2577 -4915
rect -185 -4970 2386 -4932
rect 2557 -4970 2577 -4932
rect -185 -4983 2577 -4970
rect -185 -5031 -156 -4983
rect -287 -5049 -156 -5031
rect 688 -5191 890 -5159
rect 688 -5309 724 -5191
rect 853 -5309 890 -5191
rect 688 -5339 890 -5309
rect 2233 -5308 2337 -5293
rect 2233 -5373 2249 -5308
rect 2318 -5373 2337 -5308
rect 5192 -5358 5218 -3932
rect 5945 -5306 6161 -5278
rect 2233 -5386 2337 -5373
rect 2294 -5488 2337 -5386
rect 2742 -5406 2957 -5392
rect 2742 -5442 2753 -5406
rect 2937 -5442 2957 -5406
rect 2742 -5454 2957 -5442
rect 4954 -5438 5184 -5409
rect 2294 -5514 3963 -5488
rect 2787 -5560 2988 -5553
rect 2787 -5596 2796 -5560
rect 2980 -5596 2988 -5560
rect 4954 -5555 4981 -5438
rect 5159 -5555 5184 -5438
rect 4954 -5586 5184 -5555
rect 5945 -5558 5979 -5306
rect 6123 -5558 6161 -5306
rect 5945 -5594 6161 -5558
rect 6849 -5304 7100 -5277
rect 6849 -5585 6873 -5304
rect 7061 -5585 7100 -5304
rect 2787 -5602 2988 -5596
rect 6849 -5602 7100 -5585
<< via2 >>
rect 703 1796 826 1860
rect 2791 1876 2977 1913
rect 4764 1859 5149 1912
rect 2767 1696 2953 1733
rect 4998 1735 5137 1821
rect -1456 1533 -479 1638
rect -272 1144 -226 1323
rect 2383 1309 2429 1488
rect -610 594 -532 705
rect 98 -103 397 94
rect 2046 -83 2221 91
rect 5724 1399 5786 1459
rect 2578 529 2621 751
rect 5653 753 5720 814
rect 5611 -52 5768 1
rect -268 -1350 -222 -1171
rect -1398 -1614 -1306 -1421
rect 2391 -1498 2437 -1319
rect 2581 -772 2624 -550
rect 5523 -690 5609 -609
rect 5459 -1511 5571 -1455
rect 5571 -1511 5584 -1455
rect 2754 -1739 2933 -1698
rect 709 -1908 824 -1800
rect 4972 -1940 5156 -1756
rect 2757 -2014 2936 -1973
rect -271 -2564 -225 -2385
rect 2384 -2398 2430 -2219
rect -1373 -3173 -1301 -2983
rect 67 -3810 366 -3613
rect 2035 -3767 2210 -3593
rect 2579 -3174 2622 -2952
rect 5563 -2136 5611 -2085
rect 5662 -2940 5729 -2938
rect 5662 -3000 5727 -2940
rect 5727 -3000 5729 -2940
rect 5662 -3001 5729 -3000
rect 7332 -3279 7573 -3277
rect 7332 -3315 7573 -3279
rect -268 -5031 -185 -4834
rect 2390 -4969 2548 -4933
rect 724 -5309 853 -5191
rect 2753 -5442 2937 -5406
rect 2796 -5596 2980 -5560
rect 4981 -5555 5159 -5438
rect 5979 -5558 6123 -5306
rect 6873 -5585 7061 -5304
<< metal3 >>
rect -22 1690 491 1950
rect 686 1860 847 1950
rect 686 1796 703 1860
rect 826 1796 847 1860
rect 686 1778 847 1796
rect -1483 1638 491 1690
rect -1483 1533 -1456 1638
rect -479 1533 491 1638
rect -1483 1509 491 1533
rect -287 1323 -206 1353
rect -287 1144 -272 1323
rect -226 1144 -206 1323
rect -633 705 -513 720
rect -633 594 -610 705
rect -532 594 -513 705
rect -633 578 -513 594
rect -1426 -720 -1273 -709
rect -1426 -770 -1420 -720
rect -1285 -770 -1273 -720
rect -1426 -1421 -1273 -770
rect -1426 -1614 -1398 -1421
rect -1306 -1614 -1273 -1421
rect -1426 -1638 -1273 -1614
rect -287 -1171 -206 1144
rect -287 -1350 -268 -1171
rect -222 -1350 -206 -1171
rect -287 -2385 -206 -1350
rect -287 -2564 -271 -2385
rect -225 -2564 -206 -2385
rect -1402 -2981 -1274 -2966
rect -1402 -3179 -1383 -2981
rect -1291 -3179 -1274 -2981
rect -1402 -3200 -1274 -3179
rect -287 -4816 -206 -2564
rect -22 94 491 1509
rect -22 -103 98 94
rect 397 -103 491 94
rect -22 -3613 491 -103
rect -22 -3810 67 -3613
rect 366 -3810 491 -3613
rect -287 -4834 -156 -4816
rect -287 -5031 -268 -4834
rect -185 -5031 -156 -4834
rect -287 -5049 -156 -5031
rect -287 -5622 -206 -5049
rect -22 -5621 491 -3810
rect 687 -1800 847 1778
rect 687 -1908 709 -1800
rect 824 -1908 847 -1800
rect 687 -5159 847 -1908
rect 1947 91 2307 1950
rect 2722 1913 3059 1950
rect 2722 1876 2791 1913
rect 2977 1876 3059 1913
rect 2722 1733 3059 1876
rect 2722 1696 2767 1733
rect 2953 1696 3059 1733
rect 1947 -83 2046 91
rect 2221 -83 2307 91
rect 1947 -3593 2307 -83
rect 1947 -3767 2035 -3593
rect 2210 -3767 2307 -3593
rect 687 -5191 890 -5159
rect 687 -5309 724 -5191
rect 853 -5309 890 -5191
rect 687 -5337 890 -5309
rect 688 -5339 890 -5337
rect 1947 -5621 2307 -3767
rect 2370 1488 2449 1542
rect 2370 1309 2383 1488
rect 2429 1309 2449 1488
rect 2370 -1307 2449 1309
rect 2568 751 2632 759
rect 2568 529 2578 751
rect 2621 529 2632 751
rect 2568 521 2632 529
rect 2571 -550 2635 -542
rect 2571 -772 2581 -550
rect 2624 -772 2635 -550
rect 2571 -780 2635 -772
rect 2370 -1319 2452 -1307
rect 2370 -1498 2391 -1319
rect 2437 -1498 2452 -1319
rect 2370 -1510 2452 -1498
rect 2370 -2219 2449 -1510
rect 2370 -2398 2384 -2219
rect 2430 -2398 2449 -2219
rect 2370 -4915 2449 -2398
rect 2722 -1698 3059 1696
rect 2722 -1739 2754 -1698
rect 2933 -1739 3059 -1698
rect 2722 -1973 3059 -1739
rect 2722 -2014 2757 -1973
rect 2936 -2014 3059 -1973
rect 2569 -2952 2633 -2944
rect 2569 -3174 2579 -2952
rect 2622 -3174 2633 -2952
rect 2569 -3182 2633 -3174
rect 2370 -4933 2577 -4915
rect 2370 -4969 2390 -4933
rect 2548 -4969 2577 -4933
rect 2370 -4983 2577 -4969
rect 2722 -5406 3059 -2014
rect 2722 -5442 2753 -5406
rect 2937 -5442 3059 -5406
rect 2722 -5560 3059 -5442
rect 2722 -5596 2796 -5560
rect 2980 -5596 3059 -5560
rect 2722 -5621 3059 -5596
rect 4718 1912 5231 1950
rect 4718 1859 4764 1912
rect 5149 1859 5231 1912
rect 4718 1821 5231 1859
rect 4718 1735 4998 1821
rect 5137 1735 5231 1821
rect 4718 -1756 5231 1735
rect 4718 -1940 4972 -1756
rect 5156 -1940 5231 -1756
rect 4718 -5438 5231 -1940
rect 5328 -2932 5359 1950
rect 5389 -2097 5420 1950
rect 5451 -1451 5482 1950
rect 5513 -598 5544 1950
rect 5576 5 5607 1950
rect 5638 828 5669 1950
rect 5701 1476 5732 1950
rect 5701 1459 5813 1476
rect 5701 1399 5724 1459
rect 5786 1399 5813 1459
rect 5701 1379 5813 1399
rect 5638 814 5736 828
rect 5638 753 5653 814
rect 5720 753 5736 814
rect 5638 741 5736 753
rect 5576 1 5773 5
rect 5576 -52 5611 1
rect 5768 -52 5773 1
rect 5576 -56 5773 -52
rect 5512 -609 5623 -598
rect 5512 -690 5523 -609
rect 5609 -690 5623 -609
rect 5512 -700 5623 -690
rect 5451 -1455 5590 -1451
rect 5451 -1511 5459 -1455
rect 5584 -1511 5590 -1455
rect 5451 -1517 5590 -1511
rect 5549 -2085 5624 -2071
rect 5549 -2097 5563 -2085
rect 5389 -2132 5563 -2097
rect 5549 -2136 5563 -2132
rect 5611 -2136 5624 -2085
rect 5549 -2153 5624 -2136
rect 5649 -2932 5745 -2926
rect 5328 -2938 5745 -2932
rect 5328 -2962 5662 -2938
rect 5649 -3001 5662 -2962
rect 5729 -3001 5745 -2938
rect 5649 -3014 5745 -3001
rect 4718 -5555 4981 -5438
rect 5159 -5555 5231 -5438
rect 4718 -5621 5231 -5555
rect 5919 -5306 6179 -3242
rect 5919 -5558 5979 -5306
rect 6123 -5558 6179 -5306
rect 5919 -5620 6179 -5558
rect 6826 -5304 7121 -3241
rect 6826 -5585 6873 -5304
rect 7061 -5585 7121 -5304
rect 6826 -5620 7121 -5585
rect 7318 -3277 7592 -3216
rect 7318 -3315 7332 -3277
rect 7573 -3315 7592 -3277
rect 7318 -5620 7592 -3315
<< via3 >>
rect -610 594 -532 704
rect -1420 -770 -1285 -720
rect -1383 -2983 -1291 -2981
rect -1383 -3173 -1373 -2983
rect -1373 -3173 -1301 -2983
rect -1301 -3173 -1291 -2983
rect -1383 -3179 -1291 -3173
rect 2578 529 2621 751
rect 2581 -772 2624 -550
rect 2579 -3174 2622 -2952
<< metal4 >>
rect 2568 751 2632 759
rect -632 704 -513 720
rect -632 594 -610 704
rect -532 681 -513 704
rect 2568 681 2578 751
rect -532 606 2578 681
rect -532 594 -513 606
rect -632 578 -513 594
rect 2568 529 2578 606
rect 2621 529 2632 751
rect 2568 521 2632 529
rect 2571 -550 2635 -542
rect 2571 -709 2581 -550
rect -1426 -720 2581 -709
rect -1426 -770 -1420 -720
rect -1285 -770 2581 -720
rect -1426 -772 2581 -770
rect 2624 -772 2635 -550
rect -1426 -780 2635 -772
rect 2569 -2952 2633 -2944
rect -1402 -2981 -1273 -2964
rect -1402 -3179 -1383 -2981
rect -1291 -3019 -1273 -2981
rect 2569 -3019 2579 -2952
rect -1291 -3104 2579 -3019
rect -1291 -3179 -1273 -3104
rect -1402 -3199 -1273 -3179
rect 2569 -3174 2579 -3104
rect 2622 -3174 2633 -2952
rect 2569 -3182 2633 -3174
use comp_p  comp_p_0
timestamp 1711855675
transform 1 0 1479 0 1 -736
box -1501 731 1060 2583
use comp_p  comp_p_1
timestamp 1711855675
transform 1 0 4171 0 1 -736
box -1501 731 1060 2583
use comp_p  comp_p_2
timestamp 1711855675
transform 1 0 1479 0 -1 728
box -1501 731 1060 2583
use comp_p  comp_p_3
timestamp 1711855675
transform 1 0 4171 0 -1 728
box -1501 731 1060 2583
use comp_p  comp_p_4
timestamp 1711855675
transform 1 0 1479 0 1 -4438
box -1501 731 1060 2583
use comp_p  comp_p_5
timestamp 1711855675
transform 1 0 4171 0 1 -4438
box -1501 731 1060 2583
use comp_p  comp_p_6
timestamp 1711855675
transform 1 0 4171 0 -1 -2974
box -1501 731 1060 2583
use res_ladder_vref  res_ladder_vref_0
timestamp 1762308519
transform 1 0 -2084 0 -1 -429
box 549 -1953 1704 4960
use tmux_7therm_to_3bin  tmux_7therm_to_3bin_0
timestamp 1762392494
transform 1 0 5810 0 1 1117
box -21 -4373 1875 730
use vbias_generation  vbias_generation_0
timestamp 1762372802
transform -1 0 2209 0 -1 -3359
box -142 481 1140 2133
<< labels >>
rlabel metal3 -287 -5622 -206 -4410 1 vin
port 0 n
rlabel metal1 -1535 -5389 -380 -5344 1 vref
port 1 n
rlabel metal1 7634 1408 7680 1448 1 dout0
port 2 n
rlabel metal1 7634 788 7680 828 1 dout1
port 3 n
rlabel metal1 7634 -50 7680 -10 1 dout2
port 4 n
rlabel metal3 5701 1459 5732 1950 1 d0
port 5 n
rlabel metal3 5638 814 5669 1950 1 d1
port 6 n
rlabel metal3 5576 -56 5607 1950 1 d2
port 7 n
rlabel metal3 5513 -662 5544 1950 1 d3
port 8 n
rlabel metal3 5451 -1455 5482 1950 1 d4
port 9 n
rlabel metal3 5389 -2132 5420 1950 1 d5
port 10 n
rlabel metal3 5328 -2962 5359 1950 1 d6
port 11 n
rlabel metal3 2722 1913 3059 1950 1 vdd
port 12 n
rlabel metal3 -22 94 491 1950 1 vss
port 13 n
<< end >>
