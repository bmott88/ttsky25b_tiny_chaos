* NGSPICE file created from flashADC_3bit_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9 B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_1p41 l=7
C0 R1 R2 0.01325f
C1 R2 B 0.82332f
C2 R1 B 0.82332f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ELBHUY B D S G
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 D S 0.27388f
C1 S G 0.11229f
C2 D G 0.11229f
C3 S B 0.59197f
C4 D B 0.59197f
C5 G B 0.75059f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_VTBKAA B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 S D 0.54671f
C1 S G 0.21915f
C2 G D 0.21915f
C3 S B 0.634f
C4 D B 0.634f
C5 G B 0.43443f
C6 S VSUBS 0.51455f
C7 D VSUBS 0.51455f
C8 G VSUBS 0.36418f
C9 B VSUBS 5.72384f
.ends

.subckt vbias_generation bias_n vdd XR_bias_2/R2 XR_bias_4/R1 XR_bias_3/R2 bias_p
+ vss
XXR_bias_1 vss XR_bias_2/R2 bias_p sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_2 vss XR_bias_3/R2 XR_bias_2/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_3 vss XR_bias_4/R1 XR_bias_3/R2 sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXR_bias_4 vss XR_bias_4/R1 bias_n sky130_fd_pr__res_xhigh_po_1p41_UKZ7C9
XXMn_bias vss bias_n vss bias_n sky130_fd_pr__nfet_01v8_lvt_ELBHUY
XXMp_bias vdd bias_p vdd bias_p vss sky130_fd_pr__pfet_01v8_lvt_VTBKAA
C0 vdd XR_bias_2/R2 0.01866f
C1 bias_p vdd 0.22745f
C2 XR_bias_3/R2 XR_bias_2/R2 0
C3 bias_p XR_bias_2/R2 0.05112f
C4 bias_n XR_bias_3/R2 0.06908f
C5 XR_bias_3/R2 bias_p 0.06932f
C6 XR_bias_2/R2 XR_bias_4/R1 0.06887f
C7 bias_n XR_bias_4/R1 0
C8 XR_bias_3/R2 XR_bias_4/R1 0
C9 bias_p XR_bias_4/R1 0
C10 vdd vss 6.78775f
C11 bias_n vss 2.48381f
C12 XR_bias_4/R1 vss 1.63605f
C13 XR_bias_3/R2 vss 1.57785f
C14 XR_bias_2/R2 vss 1.57097f
C15 bias_p vss 1.64123f
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_JT48NU B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_5p73 l=5.73
C0 R2 R1 0.06813f
C1 R2 B 1.74197f
C2 R1 B 1.74197f
.ends

.subckt res_ladder_vref ref2 ref5 ref6 vref ref3 ref1 ref0 ref4 vss
XXR1 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR2 vss ref6 vref sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR10 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR3 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR4 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR5 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR6 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR7 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR8 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_5p73_JT48NU
XXR9 vss ref0 vss sky130_fd_pr__res_xhigh_po_5p73_JT48NU
C0 ref3 ref5 0.06887f
C1 ref2 ref3 0
C2 ref2 ref1 0
C3 ref6 ref5 0
C4 ref1 ref0 0
C5 ref3 ref4 0
C6 ref2 ref0 0.06887f
C7 vref ref5 0.06887f
C8 vref ref6 0.16095f
C9 ref5 ref4 0
C10 ref6 ref4 0.06887f
C11 ref2 ref4 0.06887f
C12 ref1 ref3 0.06887f
C13 ref1 vss 3.4889f
C14 ref2 vss 3.42003f
C15 ref3 vss 3.42003f
C16 ref4 vss 3.42003f
C17 ref5 vss 3.42003f
C18 ref6 vss 5.161f
C19 ref0 vss 5.32418f
C20 vref vss 4.57377f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MMMA4V a_n260_n698# a_100_n500# a_n158_n500# a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n698# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
C0 a_n158_n500# a_100_n500# 0.27388f
C1 a_n158_n500# a_n100_n588# 0.11229f
C2 a_n100_n588# a_100_n500# 0.11229f
C3 a_100_n500# a_n260_n698# 0.5905f
C4 a_n158_n500# a_n260_n698# 0.5905f
C5 a_n100_n588# a_n260_n698# 0.7183f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_5VNMZ8 a_n100_n897# a_100_n800# w_n296_n1019#
+ a_n158_n800# VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 a_n100_n897# a_n158_n800# 0.17641f
C1 a_n100_n897# a_100_n800# 0.17641f
C2 a_100_n800# a_n158_n800# 0.43758f
C3 a_n100_n897# w_n296_n1019# 0.43443f
C4 w_n296_n1019# a_n158_n800# 0.51205f
C5 a_100_n800# w_n296_n1019# 0.51205f
C6 a_100_n800# VSUBS 0.41369f
C7 a_n158_n800# VSUBS 0.41369f
C8 a_n100_n897# VSUBS 0.36418f
C9 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_n158_n400# a_100_n400# 0.21931f
C1 a_n158_n400# a_n100_n488# 0.09092f
C2 a_n100_n488# a_100_n400# 0.09092f
C3 a_100_n400# a_n260_n574# 0.48057f
C4 a_n158_n400# a_n260_n574# 0.48057f
C5 a_n100_n488# a_n260_n574# 0.74751f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GUWLND a_n158_n1000# a_n100_n1097# w_n296_n1219#
+ a_100_n1000# VSUBS
X0 a_100_n1000# a_n100_n1097# a_n158_n1000# w_n296_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
C0 a_n100_n1097# a_n158_n1000# 0.21915f
C1 a_n100_n1097# a_100_n1000# 0.21915f
C2 a_100_n1000# a_n158_n1000# 0.54671f
C3 a_n100_n1097# w_n296_n1219# 0.43443f
C4 w_n296_n1219# a_n158_n1000# 0.634f
C5 a_100_n1000# w_n296_n1219# 0.634f
C6 a_100_n1000# VSUBS 0.51455f
C7 a_n158_n1000# VSUBS 0.51455f
C8 a_n100_n1097# VSUBS 0.36418f
C9 w_n296_n1219# VSUBS 5.72384f
.ends

.subckt comp_p vinp vinn vbias_p vdd tail vout latch_right out_left latch_left vss
XXMn_cs_left vss latch_right vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_out out_left vdd vdd vout vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_diode_left1 vss latch_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXMn_cs_right1 vss latch_left vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_diode_right vss latch_right vss latch_right sky130_fd_pr__nfet_01v8_lvt_AHMAL2
Xsky130_fd_pr__pfet_01v8_lvt_5VNMZ8_0 out_left vdd vdd out_left vss sky130_fd_pr__pfet_01v8_lvt_5VNMZ8
XXMn_out_left vss out_left vss latch_left sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMn_out_right vss vout vss latch_right sky130_fd_pr__nfet_01v8_lvt_MMMA4V
XXMp_tail tail vbias_p vdd vdd vss sky130_fd_pr__pfet_01v8_lvt_GUWLND
X0 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X1 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X2 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X3 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X4 tail vinp latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X5 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X6 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
X7 tail vinn latch_left vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=9.995 l=0.35
C0 vbias_p vinp 0.03011f
C1 vbias_p latch_right 0.00109f
C2 vout tail 0.00803f
C3 out_left tail 0.00652f
C4 vinp tail 2.91757f
C5 latch_right tail 8.8942f
C6 vout out_left 0.6058f
C7 latch_left vinn 1.33911f
C8 latch_left vdd 1.3971f
C9 vout vinp 0.03655f
C10 out_left vinp 0.22514f
C11 vinn vdd 2.30474f
C12 vout latch_right 0.72835f
C13 out_left latch_right 0.1431f
C14 latch_right vinp 0.51311f
C15 vbias_p latch_left 0.00103f
C16 vbias_p vinn 0.00222f
C17 vbias_p vdd 2.11961f
C18 latch_left tail 8.82993f
C19 vinn tail 0.82695f
C20 vdd tail 2.22915f
C21 vout latch_left 0.14014f
C22 out_left latch_left 0.73463f
C23 vout vinn 0.12978f
C24 out_left vinn 0.08183f
C25 vout vdd 1.62919f
C26 out_left vdd 2.99708f
C27 latch_left vinp 0.5043f
C28 latch_left latch_right 5.15792f
C29 vinn vinp 1.25697f
C30 latch_right vinn 3.53507f
C31 vdd vinp 4.26352f
C32 latch_right vdd 1.44611f
C33 vbias_p tail 0.65167f
C34 vbias_p vout 0.14426f
C35 vbias_p out_left 0.84152f
C36 vinp vss 0.4258f
C37 vinn vss 0.50566f
C38 tail vss 1.09774f
C39 vbias_p vss 0.82905f
C40 vdd vss 43.54159f
C41 vout vss 3.2381f
C42 latch_right vss 4.74799f
C43 out_left vss 3.38408f
C44 latch_left vss 5.11722f
.ends

.subckt sky130_fd_pr__pfet_01v8_A6MZLZ B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 D B 0.14266f
C1 S G 0.02934f
C2 D S 0.32105f
C3 D G 0.02934f
C4 S B 0.14266f
C5 B G 0.24043f
C6 S VSUBS 0.09023f
C7 D VSUBS 0.09023f
C8 G VSUBS 0.11914f
C9 B VSUBS 1.5811f
.ends

.subckt sky130_fd_pr__nfet_01v8_MH3LLV B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 S G 0.02545f
C1 S D 0.16211f
C2 G D 0.02545f
C3 S B 0.1317f
C4 D B 0.1317f
C5 G B 0.34289f
.ends

.subckt tmux_2to1 Y vdd XM5/G B A S vss
XXM1 vdd vdd XM5/G S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM2 vss vss XM5/G S sky130_fd_pr__nfet_01v8_MH3LLV
XXM3 vdd A Y S vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM4 vss A Y XM5/G sky130_fd_pr__nfet_01v8_MH3LLV
XXM5 vdd Y B XM5/G vss sky130_fd_pr__pfet_01v8_A6MZLZ
XXM6 vss Y B S sky130_fd_pr__nfet_01v8_MH3LLV
C0 B vdd 0.11322f
C1 XM5/G vdd 0.17343f
C2 S A 0.09932f
C3 S Y 0.13093f
C4 Y A 0.03022f
C5 S B 0.0426f
C6 Y B 0.03022f
C7 S XM5/G 0.4752f
C8 XM5/G A 0.66126f
C9 Y XM5/G 0.31571f
C10 XM5/G B 0.09611f
C11 S vdd 0.27839f
C12 vdd A 0.05809f
C13 Y vdd 0.18933f
C14 B vss 0.39578f
C15 S vss 1.22376f
C16 Y vss 0.38976f
C17 XM5/G vss 0.68597f
C18 vdd vss 4.09633f
C19 A vss 0.18036f
.ends

.subckt sky130_fd_pr__res_generic_m1_SPQYYJ R1 R2 m1_n100_n100# VSUBS
R0 R1 R2 sky130_fd_pr__res_generic_m1 w=1 l=1
C0 R2 VSUBS 0.07104f
C1 R1 VSUBS 0.07104f
C2 m1_n100_n100# VSUBS 0.10692f
.ends

.subckt inv vin vdd vout vss
XXMn vss vss vout vin sky130_fd_pr__nfet_01v8_MH3LLV
XXMp vdd vdd vout vin vss sky130_fd_pr__pfet_01v8_A6MZLZ
C0 vin vdd 0.13776f
C1 vin vout 0.12658f
C2 vdd vout 0.11998f
C3 vin vss 0.56678f
C4 vout vss 0.40687f
C5 vdd vss 1.84972f
.ends

.subckt buffer in out vdd inv_1/vin vss
Xinv_0 in vdd inv_1/vin vss inv
Xinv_1 inv_1/vin vdd out vss inv
C0 in inv_1/vin 0.01628f
C1 out vdd 0.00589f
C2 in vdd 0.01965f
C3 inv_1/vin vdd 0.16476f
C4 out inv_1/vin 0.0071f
C5 inv_1/vin vss 0.60193f
C6 out vss 0.3255f
C7 in vss 0.41789f
C8 vdd vss 3.06334f
.ends

.subckt tmux_7therm_to_3bin d0 d1 d2 d3 d4 d5 d6 q0 q1 q2 buffer_7/inv_1/vin buffer_3/inv_1/vin
+ buffer_5/out buffer_2/out buffer_4/inv_1/vin buffer_0/inv_1/vin buffer_6/out R1/R2
+ buffer_0/out buffer_5/inv_1/vin buffer_1/inv_1/vin tmux_2to1_0/XM5/G R1/R1 tmux_2to1_1/XM5/G
+ tmux_2to1_3/A tmux_2to1_2/XM5/G tmux_2to1_3/XM5/G buffer_6/inv_1/vin buffer_2/inv_1/vin
+ R1/m1_n100_n100# buffer_1/out buffer_8/in vdd vss buffer_7/in buffer_4/out
Xtmux_2to1_1 buffer_8/in vdd tmux_2to1_1/XM5/G buffer_5/out buffer_1/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_2 tmux_2to1_3/B vdd tmux_2to1_2/XM5/G buffer_6/out buffer_2/out R1/R1 vss
+ tmux_2to1
Xtmux_2to1_3 buffer_7/in vdd tmux_2to1_3/XM5/G tmux_2to1_3/B tmux_2to1_3/A buffer_8/in
+ vss tmux_2to1
XR1 R1/R1 R1/R2 R1/m1_n100_n100# vss sky130_fd_pr__res_generic_m1_SPQYYJ
Xbuffer_0 d0 buffer_0/out vdd buffer_0/inv_1/vin vss buffer
Xbuffer_1 d1 buffer_1/out vdd buffer_1/inv_1/vin vss buffer
Xbuffer_2 d2 buffer_2/out vdd buffer_2/inv_1/vin vss buffer
Xbuffer_3 d3 R1/R2 vdd buffer_3/inv_1/vin vss buffer
Xbuffer_4 d4 buffer_4/out vdd buffer_4/inv_1/vin vss buffer
Xbuffer_5 d5 buffer_5/out vdd buffer_5/inv_1/vin vss buffer
Xbuffer_6 d6 buffer_6/out vdd buffer_6/inv_1/vin vss buffer
Xbuffer_7 buffer_7/in q0 vdd buffer_7/inv_1/vin vss buffer
Xbuffer_8 buffer_8/in q1 vdd buffer_8/inv_1/vin vss buffer
Xbuffer_9 R1/R1 q2 vdd buffer_9/inv_1/vin vss buffer
Xtmux_2to1_0 tmux_2to1_3/A vdd tmux_2to1_0/XM5/G buffer_4/out buffer_0/out R1/R1 vss
+ tmux_2to1
C0 vdd R1/m1_n100_n100# 0.01544f
C1 tmux_2to1_3/A R1/R1 0.0222f
C2 buffer_4/out buffer_8/in 0.18314f
C3 vdd buffer_8/in 0.52301f
C4 R1/m1_n100_n100# R1/R2 0.0386f
C5 tmux_2to1_3/XM5/G tmux_2to1_3/B 0.0457f
C6 buffer_1/inv_1/vin R1/R1 0.02062f
C7 tmux_2to1_1/XM5/G buffer_4/out 0.02598f
C8 buffer_2/inv_1/vin tmux_2to1_3/B 0
C9 tmux_2to1_1/XM5/G vdd 0.04059f
C10 buffer_7/in tmux_2to1_3/XM5/G 0.01403f
C11 buffer_9/inv_1/vin buffer_8/inv_1/vin 0.00438f
C12 tmux_2to1_1/XM5/G tmux_2to1_2/XM5/G 0.00433f
C13 buffer_8/in buffer_1/out 0.06403f
C14 buffer_6/out buffer_3/inv_1/vin 0
C15 buffer_4/out buffer_3/inv_1/vin 0
C16 vdd buffer_3/inv_1/vin 0.32836f
C17 q2 R1/R1 0
C18 tmux_2to1_1/XM5/G buffer_1/out 0.18587f
C19 buffer_5/inv_1/vin buffer_5/out 0.00827f
C20 buffer_5/inv_1/vin buffer_4/inv_1/vin 0.00435f
C21 buffer_5/out buffer_8/inv_1/vin 0
C22 buffer_9/inv_1/vin R1/R1 0.00349f
C23 buffer_4/out tmux_2to1_3/XM5/G 0.04713f
C24 vdd tmux_2to1_3/XM5/G 0.0495f
C25 buffer_6/out d6 0.00132f
C26 tmux_2to1_1/XM5/G buffer_8/in 0.12457f
C27 d1 d2 0.00438f
C28 buffer_2/out R1/R1 0.2789f
C29 vdd d6 0.07265f
C30 vdd buffer_2/inv_1/vin 0.32649f
C31 R1/m1_n100_n100# buffer_3/inv_1/vin 0.00103f
C32 buffer_7/in q0 0
C33 buffer_8/inv_1/vin tmux_2to1_3/B 0.00974f
C34 buffer_6/out buffer_6/inv_1/vin 0.00786f
C35 vdd buffer_6/inv_1/vin 0.32835f
C36 R1/R1 d2 0.00119f
C37 buffer_7/in buffer_8/inv_1/vin 0
C38 tmux_2to1_3/A buffer_5/out 0.00456f
C39 tmux_2to1_3/XM5/G buffer_1/out 0
C40 buffer_5/out R1/R1 0.55887f
C41 tmux_2to1_3/A tmux_2to1_0/XM5/G 0.08101f
C42 tmux_2to1_0/XM5/G R1/R1 0.0674f
C43 q1 tmux_2to1_3/B 0
C44 tmux_2to1_3/A tmux_2to1_3/B 0.0101f
C45 buffer_7/in q1 0
C46 tmux_2to1_3/XM5/G buffer_8/in 0.34642f
C47 R1/R1 tmux_2to1_3/B 0.24354f
C48 buffer_0/inv_1/vin tmux_2to1_3/A 0
C49 buffer_7/in tmux_2to1_3/A 0.38438f
C50 vdd q0 0.01294f
C51 buffer_0/inv_1/vin R1/R1 0.01886f
C52 buffer_6/out buffer_5/inv_1/vin 0
C53 buffer_7/in R1/R1 0.00295f
C54 vdd buffer_5/inv_1/vin 0.32846f
C55 vdd buffer_8/inv_1/vin 0.02538f
C56 buffer_0/inv_1/vin buffer_1/inv_1/vin 0.00435f
C57 d5 buffer_5/out 0.00133f
C58 buffer_2/out d2 0
C59 q2 tmux_2to1_3/B 0
C60 buffer_2/inv_1/vin buffer_3/inv_1/vin 0.00435f
C61 tmux_2to1_3/A buffer_0/out 0.05826f
C62 vdd d1 0.07265f
C63 buffer_2/out buffer_5/out 0.05213f
C64 vdd q1 0.01294f
C65 R1/R1 buffer_0/out 0.11396f
C66 tmux_2to1_3/A buffer_4/out 0.6033f
C67 vdd tmux_2to1_3/A 0.31099f
C68 buffer_7/inv_1/vin buffer_8/inv_1/vin 0.00435f
C69 R1/R1 d3 0
C70 buffer_6/out R1/R1 0.20693f
C71 buffer_4/out R1/R1 0.26729f
C72 vdd R1/R1 2.20161f
C73 d0 d1 0.00435f
C74 buffer_9/inv_1/vin tmux_2to1_3/B 0.00176f
C75 tmux_2to1_2/XM5/G R1/R1 0.26532f
C76 buffer_8/in buffer_8/inv_1/vin 0.01384f
C77 R1/R1 R1/R2 0.03366f
C78 buffer_2/out tmux_2to1_3/B 0.04026f
C79 vdd buffer_1/inv_1/vin 0.32649f
C80 d1 buffer_1/out 0.00148f
C81 d0 tmux_2to1_3/A 0
C82 buffer_5/out buffer_4/inv_1/vin 0
C83 d0 R1/R1 0
C84 tmux_2to1_3/A buffer_1/out 0
C85 d5 d4 0.00435f
C86 d2 tmux_2to1_3/B 0
C87 R1/R1 buffer_1/out 0.22519f
C88 vdd q2 0.01294f
C89 buffer_7/inv_1/vin tmux_2to1_3/A 0
C90 d1 buffer_8/in 0
C91 buffer_5/out tmux_2to1_3/B 0.16421f
C92 buffer_1/inv_1/vin buffer_1/out 0.0086f
C93 q1 buffer_8/in 0
C94 buffer_7/in buffer_5/out 0.00264f
C95 tmux_2to1_3/A buffer_8/in 0.1382f
C96 vdd d5 0.07265f
C97 R1/m1_n100_n100# R1/R1 0.04565f
C98 R1/R1 buffer_8/in 0.07792f
C99 buffer_0/inv_1/vin tmux_2to1_0/XM5/G 0
C100 buffer_7/in tmux_2to1_0/XM5/G 0.00597f
C101 buffer_6/out buffer_9/inv_1/vin 0.00222f
C102 vdd buffer_9/inv_1/vin 0.03021f
C103 buffer_1/inv_1/vin buffer_8/in 0
C104 tmux_2to1_1/XM5/G tmux_2to1_3/A 0
C105 buffer_2/out buffer_4/out 0.0018f
C106 buffer_2/out buffer_6/out 0.01539f
C107 buffer_2/out vdd 0.64599f
C108 tmux_2to1_1/XM5/G R1/R1 0.13419f
C109 buffer_7/in tmux_2to1_3/B 0.20877f
C110 buffer_2/out tmux_2to1_2/XM5/G 0.14365f
C111 d2 d3 0.00435f
C112 vdd d2 0.07265f
C113 R1/R1 buffer_3/inv_1/vin 0.00894f
C114 buffer_5/inv_1/vin buffer_6/inv_1/vin 0.00438f
C115 buffer_6/out buffer_5/out 0.48724f
C116 buffer_4/out buffer_5/out 1.95899f
C117 vdd buffer_5/out 1.92707f
C118 buffer_6/out buffer_4/inv_1/vin 0
C119 tmux_2to1_0/XM5/G buffer_0/out 0.18135f
C120 buffer_4/out buffer_4/inv_1/vin 0.00786f
C121 vdd buffer_4/inv_1/vin 0.32846f
C122 tmux_2to1_2/XM5/G buffer_5/out 0.09828f
C123 tmux_2to1_0/XM5/G buffer_4/out 0.02654f
C124 buffer_5/out R1/R2 0.01212f
C125 vdd tmux_2to1_0/XM5/G 0.05854f
C126 tmux_2to1_3/A tmux_2to1_3/XM5/G 0.04146f
C127 buffer_0/inv_1/vin buffer_0/out 0.00873f
C128 buffer_6/out tmux_2to1_3/B 0.18281f
C129 buffer_7/in buffer_0/out 0
C130 buffer_4/out tmux_2to1_3/B 0.27938f
C131 tmux_2to1_3/XM5/G R1/R1 0
C132 vdd tmux_2to1_3/B 1.44834f
C133 buffer_5/out buffer_1/out 0.05669f
C134 d0 tmux_2to1_0/XM5/G 0
C135 buffer_2/inv_1/vin R1/R1 0.02182f
C136 buffer_7/in buffer_4/out 0.04488f
C137 buffer_0/inv_1/vin vdd 0.32203f
C138 buffer_7/in vdd 0.23539f
C139 tmux_2to1_2/XM5/G tmux_2to1_3/B 0.03416f
C140 buffer_2/inv_1/vin buffer_1/inv_1/vin 0.00438f
C141 R1/m1_n100_n100# buffer_5/out 0.01185f
C142 buffer_5/out buffer_8/in 0.33947f
C143 buffer_1/out tmux_2to1_3/B 0
C144 d4 d3 0.00438f
C145 buffer_4/out d4 0.00132f
C146 vdd d4 0.07265f
C147 buffer_7/in buffer_1/out 0
C148 tmux_2to1_1/XM5/G buffer_5/out 0.02579f
C149 buffer_4/out buffer_0/out 0.0414f
C150 buffer_7/inv_1/vin buffer_7/in 0.00796f
C151 vdd buffer_0/out 0.83616f
C152 d6 d5 0.00438f
C153 buffer_8/in tmux_2to1_3/B 0.28179f
C154 vdd d3 0.07265f
C155 buffer_6/out buffer_4/out 1.41424f
C156 tmux_2to1_3/A q0 0
C157 buffer_6/out vdd 2.9681f
C158 tmux_2to1_1/XM5/G tmux_2to1_0/XM5/G 0.00433f
C159 vdd buffer_4/out 1.75243f
C160 buffer_5/out buffer_3/inv_1/vin 0
C161 buffer_7/in buffer_8/in 0.24628f
C162 buffer_4/inv_1/vin buffer_3/inv_1/vin 0.00438f
C163 buffer_6/out tmux_2to1_2/XM5/G 0.02333f
C164 tmux_2to1_2/XM5/G buffer_4/out 0.07683f
C165 d0 buffer_0/out 0.0015f
C166 vdd tmux_2to1_2/XM5/G 0.05427f
C167 buffer_6/out R1/R2 0.00154f
C168 buffer_4/out R1/R2 0.00232f
C169 vdd R1/R2 0.32828f
C170 tmux_2to1_1/XM5/G tmux_2to1_3/B 0
C171 buffer_2/out buffer_2/inv_1/vin 0.00356f
C172 d0 vdd 0.0683f
C173 buffer_7/in tmux_2to1_1/XM5/G 0
C174 buffer_4/out buffer_1/out 0.00456f
C175 vdd buffer_1/out 0.83708f
C176 buffer_7/inv_1/vin buffer_4/out 0.00238f
C177 tmux_2to1_3/XM5/G buffer_5/out 0.01262f
C178 buffer_7/inv_1/vin vdd 0.02382f
C179 d1 R1/R1 0
C180 buffer_6/out R1/m1_n100_n100# 0
C181 R1/m1_n100_n100# buffer_4/out 0.00131f
C182 tmux_2to1_3/A vss 0.7137f
C183 tmux_2to1_0/XM5/G vss 0.55203f
C184 buffer_9/inv_1/vin vss 0.83718f
C185 q2 vss 0.40182f
C186 buffer_8/inv_1/vin vss 0.83586f
C187 q1 vss 0.40182f
C188 buffer_7/inv_1/vin vss 0.83588f
C189 q0 vss 0.40182f
C190 buffer_6/inv_1/vin vss 0.54713f
C191 buffer_6/out vss 1.02817f
C192 d6 vss 0.42023f
C193 buffer_5/inv_1/vin vss 0.54811f
C194 buffer_5/out vss 1.10288f
C195 d5 vss 0.41693f
C196 vdd vss 81.55533f
C197 buffer_4/inv_1/vin vss 0.54811f
C198 buffer_4/out vss 1.13783f
C199 d4 vss 0.41693f
C200 buffer_3/inv_1/vin vss 0.54811f
C201 R1/R2 vss 0.24595f
C202 d3 vss 0.41694f
C203 buffer_2/inv_1/vin vss 0.55981f
C204 buffer_2/out vss 0.38944f
C205 d2 vss 0.41693f
C206 buffer_1/inv_1/vin vss 0.55981f
C207 buffer_1/out vss 0.403f
C208 d1 vss 0.41693f
C209 buffer_0/inv_1/vin vss 0.55981f
C210 buffer_0/out vss 0.40723f
C211 d0 vss 0.42457f
C212 R1/m1_n100_n100# vss 0.11104f
C213 buffer_8/in vss 1.94693f
C214 buffer_7/in vss 1.30882f
C215 tmux_2to1_3/XM5/G vss 0.55181f
C216 R1/R1 vss 4.97016f
C217 tmux_2to1_3/B vss 1.00035f
C218 tmux_2to1_2/XM5/G vss 0.54992f
C219 tmux_2to1_1/XM5/G vss 0.55178f
.ends

.subckt flashADC_3bit_extracted vin vref dout0 dout1 dout2 d0 d1 d2 d3 d4 d5 d6 vdd
+ vss
Xvbias_generation_0 vbias_generation_0/bias_n vdd vbias_generation_0/XR_bias_2/R2
+ vbias_generation_0/XR_bias_4/R1 vbias_generation_0/XR_bias_3/R2 comp_p_6/vbias_p
+ vss vbias_generation
Xres_ladder_vref_0 comp_p_2/vinn comp_p_5/vinn comp_p_6/vinn vref comp_p_3/vinn comp_p_0/vinn
+ comp_p_1/vinn comp_p_4/vinn vss res_ladder_vref
Xcomp_p_1 vin comp_p_1/vinn comp_p_6/vbias_p vdd comp_p_1/tail d0 comp_p_1/latch_right
+ comp_p_1/out_left comp_p_1/latch_left vss comp_p
Xcomp_p_0 vin comp_p_0/vinn comp_p_6/vbias_p vdd comp_p_0/tail d1 comp_p_0/latch_right
+ comp_p_0/out_left comp_p_0/latch_left vss comp_p
Xcomp_p_2 vin comp_p_2/vinn comp_p_6/vbias_p vdd comp_p_2/tail d2 comp_p_2/latch_right
+ comp_p_2/out_left comp_p_2/latch_left vss comp_p
Xcomp_p_3 vin comp_p_3/vinn comp_p_6/vbias_p vdd comp_p_3/tail d3 comp_p_3/latch_right
+ comp_p_3/out_left comp_p_3/latch_left vss comp_p
Xcomp_p_4 vin comp_p_4/vinn comp_p_6/vbias_p vdd comp_p_4/tail d4 comp_p_4/latch_right
+ comp_p_4/out_left comp_p_4/latch_left vss comp_p
Xcomp_p_5 vin comp_p_5/vinn comp_p_6/vbias_p vdd comp_p_5/tail d5 comp_p_5/latch_right
+ comp_p_5/out_left comp_p_5/latch_left vss comp_p
Xcomp_p_6 vin comp_p_6/vinn comp_p_6/vbias_p vdd comp_p_6/tail d6 comp_p_6/latch_right
+ comp_p_6/out_left comp_p_6/latch_left vss comp_p
Xtmux_7therm_to_3bin_0 d0 d1 d2 d3 d4 d5 d6 dout0 dout1 dout2 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_3/inv_1/vin tmux_7therm_to_3bin_0/buffer_5/out tmux_7therm_to_3bin_0/buffer_2/out
+ tmux_7therm_to_3bin_0/buffer_4/inv_1/vin tmux_7therm_to_3bin_0/buffer_0/inv_1/vin
+ tmux_7therm_to_3bin_0/buffer_6/out tmux_7therm_to_3bin_0/R1/R2 tmux_7therm_to_3bin_0/buffer_0/out
+ tmux_7therm_to_3bin_0/buffer_5/inv_1/vin tmux_7therm_to_3bin_0/buffer_1/inv_1/vin
+ tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G tmux_7therm_to_3bin_0/R1/R1 tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G
+ tmux_7therm_to_3bin_0/tmux_2to1_3/A tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G
+ tmux_7therm_to_3bin_0/buffer_6/inv_1/vin tmux_7therm_to_3bin_0/buffer_2/inv_1/vin
+ tmux_7therm_to_3bin_0/R1/m1_n100_n100# tmux_7therm_to_3bin_0/buffer_1/out tmux_7therm_to_3bin_0/buffer_8/in
+ vdd vss tmux_7therm_to_3bin_0/buffer_7/in tmux_7therm_to_3bin_0/buffer_4/out tmux_7therm_to_3bin
X0 vdd comp_p_4/out_left.t2 d4 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X1 comp_p_5/latch_right.t1 comp_p_5/latch_right.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X2 vdd comp_p_6/out_left.t2 d6 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X3 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d1.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X4 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X5 comp_p_1/out_left comp_p_1/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X6 comp_p_2/tail vin.t10 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X7 comp_p_4/tail vin.t16 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X8 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X9 comp_p_2/tail vin.t9 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X10 vdd comp_p_6/vbias_p.t3 comp_p_0/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X11 comp_p_1/tail vin.t2 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X12 comp_p_4/tail vin.t19 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X13 comp_p_5/latch_right comp_p_5/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X14 d5 comp_p_5/latch_right.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X15 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X16 comp_p_0/latch_left comp_p_0/latch_right.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X17 comp_p_2/latch_right comp_p_2/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X18 comp_p_2/tail vin.t11 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X19 vdd comp_p_6/vbias_p.t5 comp_p_3/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X20 comp_p_1/tail vin.t3 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X21 vdd comp_p_2/out_left.t0 comp_p_2/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X22 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d1.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X23 vdd comp_p_0/out_left.t0 comp_p_0/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X24 comp_p_2/latch_left.t1 comp_p_2/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X25 comp_p_3/out_left comp_p_3/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X26 vdd comp_p_6/vbias_p.t6 comp_p_4/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X27 comp_p_4/tail vin.t18 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X28 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d3.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X29 comp_p_3/latch_left.t1 comp_p_3/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X30 vdd comp_p_6/vbias_p.t8 comp_p_6/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X31 comp_p_6/tail vin.t24 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X32 comp_p_0/tail vin.t6 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X33 vdd comp_p_6/out_left.t0 comp_p_6/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X34 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d2.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X35 comp_p_0/tail vin.t4 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X36 comp_p_3/tail vin.t12 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X37 vdd comp_p_4/out_left.t0 comp_p_4/out_left.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X38 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d2.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X39 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d3.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X40 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d5.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X41 comp_p_0/tail vin.t7 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X42 comp_p_5/tail vin.t21 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X43 comp_p_1/latch_right comp_p_1/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X44 comp_p_0/latch_right.t1 comp_p_0/latch_right.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X45 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d5.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X46 comp_p_0/tail vin.t5 comp_p_0/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X47 comp_p_1/latch_left.t1 comp_p_1/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X48 vdd comp_p_6/vbias_p.t2 comp_p_1/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X49 vdd comp_p_0/out_left.t2 d1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X50 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d0.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X51 comp_p_5/out_left comp_p_5/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X52 vdd comp_p_6/vbias_p.t4 comp_p_2/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X53 comp_p_3/latch_right comp_p_3/latch_left.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X54 comp_p_5/latch_left.t1 comp_p_5/latch_left.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=0 l=0
X55 comp_p_6/tail vin.t25 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X56 comp_p_5/latch_left comp_p_5/latch_right.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X57 comp_p_6/tail vin.t26 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X58 comp_p_2/tail vin.t8 comp_p_2/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X59 comp_p_4/tail vin.t17 comp_p_4/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X60 comp_p_5/tail vin.t20 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X61 d1 comp_p_0/latch_right.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X62 comp_p_3/tail vin.t13 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X63 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d0.t0 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X64 comp_p_3/tail vin.t14 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X65 vdd comp_p_6/vbias_p.t7 comp_p_5/tail vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X66 comp_p_6/tail vin.t27 comp_p_6/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X67 vdd comp_p_2/out_left.t2 d2 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=0 l=0
X68 comp_p_2/out_left comp_p_2/latch_left.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=0 l=0
X69 comp_p_1/tail vin.t0 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X70 vdd comp_p_6/vbias_p.t0 comp_p_6/vbias_p.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=0 l=0
X71 comp_p_5/tail vin.t23 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X72 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4.t1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
X73 comp_p_3/tail vin.t15 comp_p_3/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X74 comp_p_5/tail vin.t22 comp_p_5/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
X75 comp_p_1/tail vin.t1 comp_p_1/latch_right vdd sky130_fd_pr__pfet_01v8_lvt ad=2.89855 pd=20.57 as=2.89855 ps=20.57 w=0 l=0
R0 comp_p_6/vbias_p.t0 comp_p_6/vbias_p.n6 337.106
R1 comp_p_6/vbias_p comp_p_6/vbias_p.t0 332.425
R2 comp_p_6/vbias_p comp_p_6/vbias_p.t2 178.793
R3 comp_p_6/vbias_p comp_p_6/vbias_p.t8 178.793
R4 comp_p_6/vbias_p.n2 comp_p_6/vbias_p.t7 172.639
R5 comp_p_6/vbias_p.n2 comp_p_6/vbias_p.t5 172.639
R6 comp_p_6/vbias_p.n3 comp_p_6/vbias_p.t6 172.639
R7 comp_p_6/vbias_p.n3 comp_p_6/vbias_p.t4 172.639
R8 comp_p_6/vbias_p.n0 comp_p_6/vbias_p.t3 172.639
R9 comp_p_6/vbias_p comp_p_6/vbias_p.t1 23.0294
R10 comp_p_6/vbias_p.n8 comp_p_6/vbias_p 8.71581
R11 comp_p_6/vbias_p.n0 comp_p_6/vbias_p 6.78896
R12 comp_p_6/vbias_p.n7 comp_p_6/vbias_p 4.65471
R13 comp_p_6/vbias_p.n1 comp_p_6/vbias_p 3.50247
R14 comp_p_6/vbias_p.n7 comp_p_6/vbias_p 3.11545
R15 comp_p_6/vbias_p comp_p_6/vbias_p.n8 2.28805
R16 comp_p_6/vbias_p.n5 comp_p_6/vbias_p.n1 2.21866
R17 comp_p_6/vbias_p comp_p_6/vbias_p.n5 2.14383
R18 comp_p_6/vbias_p.n1 comp_p_6/vbias_p.n0 2.08314
R19 comp_p_6/vbias_p.n3 comp_p_6/vbias_p 1.28874
R20 comp_p_6/vbias_p comp_p_6/vbias_p.n2 1.15992
R21 comp_p_6/vbias_p.n6 comp_p_6/vbias_p 0.802583
R22 comp_p_6/vbias_p.n4 comp_p_6/vbias_p 0.714721
R23 comp_p_6/vbias_p.n8 comp_p_6/vbias_p.n7 0.451639
R24 comp_p_6/vbias_p.n4 comp_p_6/vbias_p.n3 0.445699
R25 comp_p_6/vbias_p.n5 comp_p_6/vbias_p.n4 0.379389
R26 comp_p_6/vbias_p.n6 comp_p_6/vbias_p 0.0564593
R27 vss.n880 vss.n879 296849
R28 vss.n878 vss.n877 15045.2
R29 vss.n877 vss.n299 11496.8
R30 vss.n62 vss.n47 10261.4
R31 vss.n62 vss.n31 10261.4
R32 vss.n117 vss.n37 10261.4
R33 vss.n111 vss.n37 10261.4
R34 vss.n902 vss.n899 8494.18
R35 vss.n923 vss.n882 8494.18
R36 vss.n923 vss.n883 8494.18
R37 vss.n880 vss.n300 8395.1
R38 vss.n907 vss.n906 7120.97
R39 vss.n906 vss.n894 7120.97
R40 vss.n912 vss.n891 7120.97
R41 vss.n912 vss.n911 7120.97
R42 vss.n918 vss.n886 7120.97
R43 vss.n918 vss.n887 7120.97
R44 vss.n74 vss.n72 6385.12
R45 vss.n74 vss.n73 6385.12
R46 vss.n67 vss.n65 6385.12
R47 vss.n67 vss.n66 6385.12
R48 vss.n80 vss.n78 6385.12
R49 vss.n80 vss.n79 6385.12
R50 vss.n57 vss.n55 6385.12
R51 vss.n57 vss.n56 6385.12
R52 vss.n95 vss.n93 6385.12
R53 vss.n95 vss.n94 6385.12
R54 vss.n89 vss.n87 6385.12
R55 vss.n89 vss.n88 6385.12
R56 vss.n106 vss.n105 6385.12
R57 vss.n106 vss.n52 6385.12
R58 vss.n100 vss.n99 6385.12
R59 vss.n100 vss.n51 6385.12
R60 vss.n113 vss.n38 6385.12
R61 vss.n113 vss.n112 6385.12
R62 vss.n283 vss.n169 5440.68
R63 vss.n947 vss.n167 5440.68
R64 vss.n214 vss.n155 5440.68
R65 vss.n160 vss.n158 5440.68
R66 vss.n808 vss.n620 5440.68
R67 vss.n745 vss.n743 5440.68
R68 vss.n806 vss.n628 5440.68
R69 vss.n251 vss.n170 5255.26
R70 vss.n945 vss.n171 5255.26
R71 vss.n958 vss.n151 5255.26
R72 vss.n956 vss.n955 5255.26
R73 vss.n664 vss.n649 5255.26
R74 vss.n783 vss.n723 5255.26
R75 vss.n701 vss.n652 5255.26
R76 vss.n714 vss.n296 5116.21
R77 vss.n714 vss.n294 5116.21
R78 vss.n926 vss.n296 5116.21
R79 vss.n926 vss.n294 5116.21
R80 vss.n879 vss.n878 4557.71
R81 vss.n225 vss.n181 4536.79
R82 vss.n268 vss.n225 4536.79
R83 vss.n273 vss.n174 4536.79
R84 vss.n940 vss.n174 4536.79
R85 vss.n237 vss.n228 4536.79
R86 vss.n228 vss.n177 4536.79
R87 vss.n966 vss.n121 4536.79
R88 vss.n121 vss.n18 4536.79
R89 vss.n126 vss.n15 4536.79
R90 vss.n134 vss.n126 4536.79
R91 vss.n968 vss.n20 4536.79
R92 vss.n981 vss.n20 4536.79
R93 vss.n713 vss.n639 4536.79
R94 vss.n793 vss.n639 4536.79
R95 vss.n660 vss.n659 4536.79
R96 vss.n684 vss.n660 4536.79
R97 vss.n788 vss.n717 4536.79
R98 vss.n788 vss.n718 4536.79
R99 vss.n769 vss.n739 4536.79
R100 vss.n769 vss.n737 4536.79
R101 vss.n686 vss.n656 4536.79
R102 vss.n688 vss.n656 4536.79
R103 vss.n790 vss.n712 4536.79
R104 vss.n790 vss.n630 4536.79
R105 vss.n246 vss.n170 4131.21
R106 vss.n245 vss.n178 4131.21
R107 vss.n282 vss.n180 4131.21
R108 vss.n240 vss.n238 4131.21
R109 vss.n241 vss.n220 4131.21
R110 vss.n945 vss.n166 4131.21
R111 vss.n234 vss.n229 4131.21
R112 vss.n275 vss.n233 4131.21
R113 vss.n182 vss.n176 4131.21
R114 vss.n938 vss.n183 4131.21
R115 vss.n213 vss.n151 4131.21
R116 vss.n137 vss.n135 4131.21
R117 vss.n139 vss.n138 4131.21
R118 vss.n16 vss.n11 4131.21
R119 vss.n983 vss.n12 4131.21
R120 vss.n955 vss.n159 4131.21
R121 vss.n133 vss.n128 4131.21
R122 vss.n970 vss.n132 4131.21
R123 vss.n127 vss.n14 4131.21
R124 vss.n157 vss.n19 4131.21
R125 vss.n649 vss.n619 4131.21
R126 vss.n670 vss.n651 4131.21
R127 vss.n794 vss.n626 4131.21
R128 vss.n669 vss.n650 4131.21
R129 vss.n638 vss.n624 4131.21
R130 vss.n726 vss.n723 4131.21
R131 vss.n758 vss.n757 4131.21
R132 vss.n760 vss.n759 4131.21
R133 vss.n732 vss.n725 4131.21
R134 vss.n766 vss.n746 4131.21
R135 vss.n701 vss.n627 4131.21
R136 vss.n703 vss.n646 4131.21
R137 vss.n642 vss.n622 4131.21
R138 vss.n696 vss.n648 4131.21
R139 vss.n707 vss.n623 4131.21
R140 vss.n575 vss.n574 4116.13
R141 vss.n246 vss.n169 3945.79
R142 vss.n250 vss.n178 3945.79
R143 vss.n245 vss.n180 3945.79
R144 vss.n242 vss.n238 3945.79
R145 vss.n241 vss.n240 3945.79
R146 vss.n947 vss.n166 3945.79
R147 vss.n269 vss.n234 3945.79
R148 vss.n275 vss.n229 3945.79
R149 vss.n176 vss.n175 3945.79
R150 vss.n938 vss.n182 3945.79
R151 vss.n214 vss.n213 3945.79
R152 vss.n140 vss.n135 3945.79
R153 vss.n139 vss.n137 3945.79
R154 vss.n152 vss.n16 3945.79
R155 vss.n983 vss.n11 3945.79
R156 vss.n160 vss.n159 3945.79
R157 vss.n133 vss.n26 3945.79
R158 vss.n970 vss.n128 3945.79
R159 vss.n21 vss.n14 3945.79
R160 vss.n127 vss.n19 3945.79
R161 vss.n808 vss.n619 3945.79
R162 vss.n677 vss.n651 3945.79
R163 vss.n670 vss.n626 3945.79
R164 vss.n661 vss.n650 3945.79
R165 vss.n669 vss.n624 3945.79
R166 vss.n743 vss.n726 3945.79
R167 vss.n757 vss.n750 3945.79
R168 vss.n760 vss.n758 3945.79
R169 vss.n732 vss.n722 3945.79
R170 vss.n766 vss.n725 3945.79
R171 vss.n806 vss.n627 3945.79
R172 vss.n703 vss.n645 3945.79
R173 vss.n646 vss.n622 3945.79
R174 vss.n658 vss.n648 3945.79
R175 vss.n696 vss.n623 3945.79
R176 vss.n52 vss.n44 3876.26
R177 vss.n94 vss.n44 3876.26
R178 vss.n79 vss.n46 3876.26
R179 vss.n73 vss.n46 3876.26
R180 vss.n66 vss.n47 3876.26
R181 vss.n72 vss.n33 3876.26
R182 vss.n65 vss.n33 3876.26
R183 vss.n65 vss.n31 3876.26
R184 vss.n73 vss.n48 3876.26
R185 vss.n66 vss.n48 3876.26
R186 vss.n55 vss.n34 3876.26
R187 vss.n78 vss.n34 3876.26
R188 vss.n78 vss.n30 3876.26
R189 vss.n72 vss.n30 3876.26
R190 vss.n88 vss.n45 3876.26
R191 vss.n56 vss.n45 3876.26
R192 vss.n56 vss.n49 3876.26
R193 vss.n79 vss.n49 3876.26
R194 vss.n93 vss.n35 3876.26
R195 vss.n87 vss.n35 3876.26
R196 vss.n87 vss.n29 3876.26
R197 vss.n55 vss.n29 3876.26
R198 vss.n94 vss.n50 3876.26
R199 vss.n88 vss.n50 3876.26
R200 vss.n99 vss.n36 3876.26
R201 vss.n105 vss.n36 3876.26
R202 vss.n105 vss.n28 3876.26
R203 vss.n93 vss.n28 3876.26
R204 vss.n112 vss.n42 3876.26
R205 vss.n51 vss.n42 3876.26
R206 vss.n109 vss.n51 3876.26
R207 vss.n109 vss.n52 3876.26
R208 vss.n117 vss.n38 3876.26
R209 vss.n38 vss.n27 3876.26
R210 vss.n99 vss.n27 3876.26
R211 vss.n112 vss.n111 3876.26
R212 vss.n250 vss.n181 3227.32
R213 vss.n268 vss.n242 3227.32
R214 vss.n239 vss.n220 3227.32
R215 vss.n273 vss.n269 3227.32
R216 vss.n237 vss.n233 3227.32
R217 vss.n940 vss.n175 3227.32
R218 vss.n183 vss.n177 3227.32
R219 vss.n966 vss.n140 3227.32
R220 vss.n138 vss.n136 3227.32
R221 vss.n152 vss.n18 3227.32
R222 vss.n968 vss.n26 3227.32
R223 vss.n134 vss.n132 3227.32
R224 vss.n981 vss.n21 3227.32
R225 vss.n157 vss.n15 3227.32
R226 vss.n677 vss.n659 3227.32
R227 vss.n794 vss.n793 3227.32
R228 vss.n684 vss.n661 3227.32
R229 vss.n713 vss.n638 3227.32
R230 vss.n750 vss.n717 3227.32
R231 vss.n759 vss.n739 3227.32
R232 vss.n722 vss.n718 3227.32
R233 vss.n746 vss.n737 3227.32
R234 vss.n686 vss.n645 3227.32
R235 vss.n712 vss.n642 3227.32
R236 vss.n688 vss.n658 3227.32
R237 vss.n707 vss.n630 3227.32
R238 vss.n880 vss.n299 2649.46
R239 vss.n879 vss.n301 2447.15
R240 vss.n361 vss.n344 2306.06
R241 vss.n347 vss.n344 2306.06
R242 vss.n361 vss.n345 2306.06
R243 vss.n347 vss.n345 2306.06
R244 vss.n371 vss.n334 2306.06
R245 vss.n363 vss.n334 2306.06
R246 vss.n371 vss.n335 2306.06
R247 vss.n363 vss.n335 2306.06
R248 vss.n473 vss.n469 2306.06
R249 vss.n473 vss.n470 2306.06
R250 vss.n483 vss.n329 2306.06
R251 vss.n330 vss.n329 2306.06
R252 vss.n435 vss.n408 2306.06
R253 vss.n450 vss.n408 2306.06
R254 vss.n435 vss.n409 2306.06
R255 vss.n450 vss.n409 2306.06
R256 vss.n422 vss.n415 2306.06
R257 vss.n432 vss.n415 2306.06
R258 vss.n422 vss.n416 2306.06
R259 vss.n432 vss.n416 2306.06
R260 vss.n352 vss.n342 2306.06
R261 vss.n354 vss.n352 2306.06
R262 vss.n353 vss.n342 2306.06
R263 vss.n354 vss.n353 2306.06
R264 vss.n340 vss.n332 2306.06
R265 vss.n365 vss.n340 2306.06
R266 vss.n341 vss.n332 2306.06
R267 vss.n365 vss.n341 2306.06
R268 vss.n475 vss.n386 2306.06
R269 vss.n475 vss.n390 2306.06
R270 vss.n481 vss.n375 2306.06
R271 vss.n375 vss.n331 2306.06
R272 vss.n447 vss.n443 2306.06
R273 vss.n447 vss.n444 2306.06
R274 vss.n466 vss.n392 2306.06
R275 vss.n466 vss.n393 2306.06
R276 vss.n437 vss.n411 2306.06
R277 vss.n441 vss.n411 2306.06
R278 vss.n437 vss.n412 2306.06
R279 vss.n441 vss.n412 2306.06
R280 vss.n424 vss.n420 2306.06
R281 vss.n420 vss.n414 2306.06
R282 vss.n425 vss.n424 2306.06
R283 vss.n425 vss.n414 2306.06
R284 vss.n868 vss.n849 2306.06
R285 vss.n849 vss.n846 2306.06
R286 vss.n868 vss.n850 2306.06
R287 vss.n850 vss.n846 2306.06
R288 vss.n848 vss.n843 2306.06
R289 vss.n870 vss.n843 2306.06
R290 vss.n848 vss.n844 2306.06
R291 vss.n870 vss.n844 2306.06
R292 vss.n856 vss.n304 2306.06
R293 vss.n861 vss.n304 2306.06
R294 vss.n860 vss.n856 2306.06
R295 vss.n861 vss.n860 2306.06
R296 vss.n528 vss.n508 2306.06
R297 vss.n517 vss.n508 2306.06
R298 vss.n528 vss.n509 2306.06
R299 vss.n517 vss.n509 2306.06
R300 vss.n594 vss.n530 2306.06
R301 vss.n598 vss.n530 2306.06
R302 vss.n594 vss.n531 2306.06
R303 vss.n598 vss.n531 2306.06
R304 vss.n579 vss.n548 2306.06
R305 vss.n577 vss.n548 2306.06
R306 vss.n589 vss.n533 2306.06
R307 vss.n589 vss.n534 2306.06
R308 vss.n561 vss.n550 2306.06
R309 vss.n573 vss.n550 2306.06
R310 vss.n561 vss.n551 2306.06
R311 vss.n573 vss.n551 2306.06
R312 vss.n564 vss.n554 2306.06
R313 vss.n557 vss.n555 2306.06
R314 vss.n564 vss.n555 2306.06
R315 vss.n515 vss.n506 2306.06
R316 vss.n519 vss.n515 2306.06
R317 vss.n516 vss.n506 2306.06
R318 vss.n519 vss.n516 2306.06
R319 vss.n592 vss.n503 2306.06
R320 vss.n600 vss.n503 2306.06
R321 vss.n592 vss.n504 2306.06
R322 vss.n600 vss.n504 2306.06
R323 vss.n831 vss.n819 2306.06
R324 vss.n833 vss.n819 2306.06
R325 vss.n831 vss.n820 2306.06
R326 vss.n833 vss.n820 2306.06
R327 vss.n829 vss.n823 2306.06
R328 vss.n823 vss.n822 2306.06
R329 vss.n829 vss.n824 2306.06
R330 vss.n824 vss.n822 2306.06
R331 vss.n875 vss.n306 2306.06
R332 vss.n875 vss.n307 2306.06
R333 vss.n858 vss.n306 2306.06
R334 vss.n858 vss.n307 2306.06
R335 vss.n881 vss.n298 2024.56
R336 vss.n282 vss.n179 1825.15
R337 vss.n209 vss.n12 1825.15
R338 vss.n702 vss.n621 1455.1
R339 vss.n807 vss.n625 1455.1
R340 vss.n326 vss.n322 1390.59
R341 vss.n326 vss.n316 1390.59
R342 vss.n323 vss.n321 1390.59
R343 vss.n323 vss.n315 1390.59
R344 vss.n378 vss.n374 1390.59
R345 vss.n378 vss.n377 1390.59
R346 vss.n388 vss.n387 1390.59
R347 vss.n389 vss.n388 1390.59
R348 vss.n402 vss.n401 1390.59
R349 vss.n401 vss.n397 1390.59
R350 vss.n403 vss.n400 1390.59
R351 vss.n403 vss.n396 1390.59
R352 vss.n544 vss.n543 1390.59
R353 vss.n543 vss.n539 1390.59
R354 vss.n545 vss.n542 1390.59
R355 vss.n545 vss.n538 1390.59
R356 vss.n702 vss.n647 1389.8
R357 vss.n807 vss.n621 1389.8
R358 vss.n907 vss.n896 1373.21
R359 vss.n911 vss.n910 1373.21
R360 vss.n910 vss.n894 1373.21
R361 vss.n902 vss.n894 1373.21
R362 vss.n915 vss.n886 1373.21
R363 vss.n915 vss.n891 1373.21
R364 vss.n908 vss.n891 1373.21
R365 vss.n908 vss.n907 1373.21
R366 vss.n886 vss.n882 1373.21
R367 vss.n887 vss.n883 1373.21
R368 vss.n889 vss.n887 1373.21
R369 vss.n911 vss.n889 1373.21
R370 vss.n242 vss.n227 1309.47
R371 vss.n250 vss.n227 1309.47
R372 vss.n240 vss.n226 1309.47
R373 vss.n245 vss.n226 1309.47
R374 vss.n251 vss.n250 1309.47
R375 vss.n247 vss.n245 1309.47
R376 vss.n247 vss.n246 1309.47
R377 vss.n281 vss.n220 1309.47
R378 vss.n282 vss.n281 1309.47
R379 vss.n283 vss.n282 1309.47
R380 vss.n175 vss.n171 1309.47
R381 vss.n184 vss.n182 1309.47
R382 vss.n184 vss.n166 1309.47
R383 vss.n183 vss.n167 1309.47
R384 vss.n233 vss.n224 1309.47
R385 vss.n224 vss.n183 1309.47
R386 vss.n279 vss.n229 1309.47
R387 vss.n279 vss.n182 1309.47
R388 vss.n269 vss.n223 1309.47
R389 vss.n223 vss.n175 1309.47
R390 vss.n213 vss.n156 1309.47
R391 vss.n156 vss.n11 1309.47
R392 vss.n958 vss.n152 1309.47
R393 vss.n155 vss.n12 1309.47
R394 vss.n152 vss.n125 1309.47
R395 vss.n140 vss.n125 1309.47
R396 vss.n122 vss.n11 1309.47
R397 vss.n137 vss.n122 1309.47
R398 vss.n124 vss.n12 1309.47
R399 vss.n138 vss.n124 1309.47
R400 vss.n159 vss.n154 1309.47
R401 vss.n154 vss.n127 1309.47
R402 vss.n956 vss.n21 1309.47
R403 vss.n158 vss.n157 1309.47
R404 vss.n976 vss.n21 1309.47
R405 vss.n976 vss.n26 1309.47
R406 vss.n974 vss.n127 1309.47
R407 vss.n974 vss.n128 1309.47
R408 vss.n157 vss.n120 1309.47
R409 vss.n132 vss.n120 1309.47
R410 vss.n708 vss.n642 1309.47
R411 vss.n708 vss.n707 1309.47
R412 vss.n668 vss.n619 1309.47
R413 vss.n669 vss.n668 1309.47
R414 vss.n664 vss.n661 1309.47
R415 vss.n638 vss.n620 1309.47
R416 vss.n678 vss.n661 1309.47
R417 vss.n678 vss.n677 1309.47
R418 vss.n671 vss.n669 1309.47
R419 vss.n671 vss.n670 1309.47
R420 vss.n795 vss.n638 1309.47
R421 vss.n795 vss.n794 1309.47
R422 vss.n783 vss.n722 1309.47
R423 vss.n780 vss.n725 1309.47
R424 vss.n780 vss.n726 1309.47
R425 vss.n746 vss.n745 1309.47
R426 vss.n759 vss.n741 1309.47
R427 vss.n746 vss.n741 1309.47
R428 vss.n758 vss.n749 1309.47
R429 vss.n749 vss.n725 1309.47
R430 vss.n754 vss.n750 1309.47
R431 vss.n754 vss.n722 1309.47
R432 vss.n658 vss.n652 1309.47
R433 vss.n697 vss.n696 1309.47
R434 vss.n697 vss.n627 1309.47
R435 vss.n707 vss.n628 1309.47
R436 vss.n695 vss.n646 1309.47
R437 vss.n696 vss.n695 1309.47
R438 vss.n657 vss.n645 1309.47
R439 vss.n658 vss.n657 1309.47
R440 vss.n209 vss.n208 1251.53
R441 vss.n687 vss.n302 1136.73
R442 vss.n687 vss.n647 1136.73
R443 vss.n792 vss.n625 1136.73
R444 vss.n792 vss.n791 1136.73
R445 vss.n469 vss.n321 915.471
R446 vss.n487 vss.n321 915.471
R447 vss.n487 vss.n322 915.471
R448 vss.n483 vss.n322 915.471
R449 vss.n470 vss.n315 915.471
R450 vss.n489 vss.n315 915.471
R451 vss.n489 vss.n316 915.471
R452 vss.n330 vss.n316 915.471
R453 vss.n387 vss.n386 915.471
R454 vss.n387 vss.n320 915.471
R455 vss.n374 vss.n320 915.471
R456 vss.n481 vss.n374 915.471
R457 vss.n390 vss.n389 915.471
R458 vss.n389 vss.n318 915.471
R459 vss.n377 vss.n318 915.471
R460 vss.n377 vss.n331 915.471
R461 vss.n443 vss.n400 915.471
R462 vss.n459 vss.n400 915.471
R463 vss.n459 vss.n402 915.471
R464 vss.n402 vss.n392 915.471
R465 vss.n444 vss.n396 915.471
R466 vss.n461 vss.n396 915.471
R467 vss.n461 vss.n397 915.471
R468 vss.n397 vss.n393 915.471
R469 vss.n579 vss.n542 915.471
R470 vss.n584 vss.n542 915.471
R471 vss.n584 vss.n544 915.471
R472 vss.n544 vss.n533 915.471
R473 vss.n577 vss.n538 915.471
R474 vss.n586 vss.n538 915.471
R475 vss.n586 vss.n539 915.471
R476 vss.n539 vss.n534 915.471
R477 vss.n881 vss.n880 859.029
R478 vss.n791 vss.n789 751.02
R479 vss.n929 vss.n928 705.364
R480 vss.n63 vss.n61 666.73
R481 vss vss.n63 666.73
R482 vss.n789 vss.n716 659.184
R483 vss.n116 vss.n39 621.553
R484 vss vss.n43 619.196
R485 vss.n928 vss.n927 599.019
R486 vss.n208 vss.n5 585
R487 vss.n208 vss.n17 585
R488 vss.n210 vss.n209 585
R489 vss.n209 vss.n13 585
R490 vss.n563 vss.n559 560.645
R491 vss.n562 vss.n549 560.645
R492 vss.n574 vss.n549 560.645
R493 vss.n578 vss.n575 560.645
R494 vss.n578 vss.n540 560.645
R495 vss.n585 vss.n540 560.645
R496 vss.n585 vss.n541 560.645
R497 vss.n541 vss.n532 560.645
R498 vss.n590 vss.n532 560.645
R499 vss.n593 vss.n505 560.645
R500 vss.n599 vss.n505 560.645
R501 vss.n529 vss.n507 560.645
R502 vss.n518 vss.n507 560.645
R503 vss.n423 vss.n413 560.645
R504 vss.n433 vss.n413 560.645
R505 vss.n436 vss.n410 560.645
R506 vss.n449 vss.n410 560.645
R507 vss.n448 vss.n442 560.645
R508 vss.n442 vss.n398 560.645
R509 vss.n460 vss.n398 560.645
R510 vss.n460 vss.n399 560.645
R511 vss.n399 vss.n391 560.645
R512 vss.n467 vss.n391 560.645
R513 vss.n474 vss.n468 560.645
R514 vss.n468 vss.n317 560.645
R515 vss.n488 vss.n317 560.645
R516 vss.n488 vss.n319 560.645
R517 vss.n482 vss.n319 560.645
R518 vss.n482 vss.n373 560.645
R519 vss.n372 vss.n333 560.645
R520 vss.n364 vss.n333 560.645
R521 vss.n362 vss.n343 560.645
R522 vss.n343 vss.n300 560.645
R523 vss.n898 vss 551.907
R524 vss.n903 vss.n898 551.907
R525 vss.n922 vss.n921 551.907
R526 vss.n716 vss.n715 550.859
R527 vss.n144 vss.n123 534.431
R528 vss.n261 vss.n222 531.552
R529 vss.n768 vss.n740 490.01
R530 vss.n768 vss.n767 490.01
R531 vss.n767 vss.n742 490.01
R532 vss.n742 vss.n298 490.01
R533 vss.n558 vss.n557 476.983
R534 vss.n905 vss.n897 462.683
R535 vss.n905 vss.n904 462.683
R536 vss.n914 vss.n913 462.683
R537 vss.n913 vss.n893 462.683
R538 vss.n919 vss.n885 462.683
R539 vss.n920 vss.n919 462.683
R540 vss.n917 vss.n888 435.882
R541 vss.n917 vss.n916 435.882
R542 vss.n916 vss.n890 435.882
R543 vss.n909 vss.n890 435.882
R544 vss.n909 vss.n895 435.882
R545 vss.n901 vss.n895 435.882
R546 vss.n900 vss.n899 424.591
R547 vss.n756 vss.n755 417.005
R548 vss.n755 vss.n724 417.005
R549 vss.n782 vss.n724 417.005
R550 vss.n782 vss.n781 417.005
R551 vss.n715 vss.n297 417.005
R552 vss.n925 vss.n297 417.005
R553 vss.n69 vss.n68 414.872
R554 vss.n68 vss.n64 414.872
R555 vss.n75 vss.n71 414.872
R556 vss.n76 vss.n75 414.872
R557 vss.n84 vss.n58 414.872
R558 vss.n60 vss.n58 414.872
R559 vss.n82 vss.n81 414.872
R560 vss.n81 vss.n77 414.872
R561 vss.n90 vss.n86 414.872
R562 vss.n91 vss.n90 414.872
R563 vss.n97 vss.n96 414.872
R564 vss.n96 vss.n92 414.872
R565 vss.n102 vss.n101 414.872
R566 vss.n101 vss.n53 414.872
R567 vss.n107 vss.n104 414.872
R568 vss.n108 vss.n107 414.872
R569 vss.n115 vss.n114 414.872
R570 vss.n114 vss.n41 414.872
R571 vss.n593 vss.n590 376.13
R572 vss.n449 vss.n448 376.13
R573 vss.n474 vss.n467 376.13
R574 vss.n373 vss.n372 376.13
R575 vss.n563 vss.n562 369.033
R576 vss.n599 vss.n529 369.033
R577 vss.n436 vss.n433 369.033
R578 vss.n364 vss.n362 369.033
R579 vss.n477 vss.n476 343.154
R580 vss.n888 vss.n881 339.783
R581 vss vss.n295 335.06
R582 vss.n118 vss.n32 320.18
R583 vss.n110 vss.n32 320.18
R584 vss.n832 vss.n821 298.207
R585 vss.n832 vss.n301 298.207
R586 vss.n869 vss.n845 298.207
R587 vss.n869 vss.n303 298.207
R588 vss.n876 vss.n305 298.207
R589 vss.n859 vss.n305 298.207
R590 vss.n711 vss.n631 294.776
R591 vss.n666 vss.n662 294.776
R592 vss.n641 vss.n640 294.776
R593 vss.n965 vss.n141 294.776
R594 vss.n267 vss.n243 294.776
R595 vss.n236 vss.n235 294.776
R596 vss.n967 vss.n22 294.776
R597 vss.n203 vss.n202 294.776
R598 vss.n272 vss.n173 294.776
R599 vss.n770 vss.n738 294.776
R600 vss.n787 vss.n719 294.776
R601 vss.n685 vss.n655 294.776
R602 vss.n504 vss.n502 292.5
R603 vss.n505 vss.n504 292.5
R604 vss.n503 vss 292.5
R605 vss.n505 vss.n503 292.5
R606 vss.n516 vss.n514 292.5
R607 vss.n516 vss.n507 292.5
R608 vss.n515 vss 292.5
R609 vss.n515 vss.n507 292.5
R610 vss.n555 vss 292.5
R611 vss.n559 vss.n555 292.5
R612 vss.n554 vss.n553 292.5
R613 vss vss.n551 292.5
R614 vss.n551 vss.n549 292.5
R615 vss.n552 vss.n550 292.5
R616 vss.n550 vss.n549 292.5
R617 vss vss.n534 292.5
R618 vss.n534 vss.n532 292.5
R619 vss vss.n586 292.5
R620 vss.n586 vss.n585 292.5
R621 vss.n577 vss 292.5
R622 vss.n578 vss.n577 292.5
R623 vss.n580 vss.n579 292.5
R624 vss.n579 vss.n578 292.5
R625 vss.n584 vss.n583 292.5
R626 vss.n585 vss.n584 292.5
R627 vss.n535 vss.n533 292.5
R628 vss.n533 vss.n532 292.5
R629 vss vss.n531 292.5
R630 vss.n531 vss.n505 292.5
R631 vss.n596 vss.n530 292.5
R632 vss.n530 vss.n505 292.5
R633 vss vss.n509 292.5
R634 vss.n509 vss.n507 292.5
R635 vss.n510 vss.n508 292.5
R636 vss.n508 vss.n507 292.5
R637 vss vss.n824 292.5
R638 vss.n824 vss.n301 292.5
R639 vss.n825 vss.n823 292.5
R640 vss.n823 vss.n821 292.5
R641 vss.n820 vss 292.5
R642 vss.n820 vss.n301 292.5
R643 vss.n819 vss.n818 292.5
R644 vss.n821 vss.n819 292.5
R645 vss.n860 vss.n854 292.5
R646 vss.n860 vss.n859 292.5
R647 vss vss.n304 292.5
R648 vss.n876 vss.n304 292.5
R649 vss.n844 vss 292.5
R650 vss.n844 vss.n303 292.5
R651 vss.n843 vss.n842 292.5
R652 vss.n845 vss.n843 292.5
R653 vss vss.n850 292.5
R654 vss.n850 vss.n303 292.5
R655 vss.n851 vss.n849 292.5
R656 vss.n849 vss.n845 292.5
R657 vss.n858 vss.n857 292.5
R658 vss.n859 vss.n858 292.5
R659 vss.n875 vss 292.5
R660 vss.n876 vss.n875 292.5
R661 vss.n426 vss.n425 292.5
R662 vss.n425 vss.n413 292.5
R663 vss.n420 vss 292.5
R664 vss.n420 vss.n413 292.5
R665 vss.n439 vss.n412 292.5
R666 vss.n412 vss.n410 292.5
R667 vss vss.n411 292.5
R668 vss.n411 vss.n410 292.5
R669 vss.n464 vss.n393 292.5
R670 vss.n393 vss.n391 292.5
R671 vss.n462 vss.n461 292.5
R672 vss.n461 vss.n460 292.5
R673 vss.n445 vss.n444 292.5
R674 vss.n444 vss.n442 292.5
R675 vss vss.n443 292.5
R676 vss.n443 vss.n442 292.5
R677 vss.n459 vss 292.5
R678 vss.n460 vss.n459 292.5
R679 vss vss.n392 292.5
R680 vss.n392 vss.n391 292.5
R681 vss.n381 vss.n331 292.5
R682 vss.n482 vss.n331 292.5
R683 vss.n383 vss.n318 292.5
R684 vss.n488 vss.n318 292.5
R685 vss.n390 vss.n385 292.5
R686 vss.n468 vss.n390 292.5
R687 vss.n386 vss 292.5
R688 vss.n468 vss.n386 292.5
R689 vss vss.n320 292.5
R690 vss.n488 vss.n320 292.5
R691 vss.n481 vss 292.5
R692 vss.n482 vss.n481 292.5
R693 vss.n341 vss.n339 292.5
R694 vss.n341 vss.n333 292.5
R695 vss.n340 vss 292.5
R696 vss.n340 vss.n333 292.5
R697 vss.n353 vss.n351 292.5
R698 vss.n353 vss.n343 292.5
R699 vss.n352 vss 292.5
R700 vss.n352 vss.n343 292.5
R701 vss vss.n416 292.5
R702 vss.n416 vss.n413 292.5
R703 vss.n417 vss.n415 292.5
R704 vss.n415 vss.n413 292.5
R705 vss.n409 vss 292.5
R706 vss.n410 vss.n409 292.5
R707 vss.n408 vss.n407 292.5
R708 vss.n410 vss.n408 292.5
R709 vss.n330 vss 292.5
R710 vss.n482 vss.n330 292.5
R711 vss vss.n489 292.5
R712 vss.n489 vss.n488 292.5
R713 vss vss.n470 292.5
R714 vss.n470 vss.n468 292.5
R715 vss.n471 vss.n469 292.5
R716 vss.n469 vss.n468 292.5
R717 vss.n487 vss.n486 292.5
R718 vss.n488 vss.n487 292.5
R719 vss.n484 vss.n483 292.5
R720 vss.n483 vss.n482 292.5
R721 vss vss.n335 292.5
R722 vss.n335 vss.n333 292.5
R723 vss.n336 vss.n334 292.5
R724 vss.n334 vss.n333 292.5
R725 vss vss.n345 292.5
R726 vss.n345 vss.n343 292.5
R727 vss.n346 vss.n344 292.5
R728 vss.n344 vss.n343 292.5
R729 vss vss.n293 285.604
R730 vss.n809 vss.n618 280.32
R731 vss.n215 vss.n212 280.32
R732 vss.n285 vss.n284 280.32
R733 vss.n197 vss.n161 280.32
R734 vss.n948 vss.n165 280.32
R735 vss.n744 vss.n728 280.32
R736 vss.n805 vss.n804 280.32
R737 vss.n663 vss.n617 268.425
R738 vss.n675 vss.n674 268.425
R739 vss.n673 vss.n637 268.425
R740 vss.n148 vss.n147 268.425
R741 vss.n146 vss.n145 268.425
R742 vss.n207 vss.n150 268.425
R743 vss.n249 vss.n218 268.425
R744 vss.n265 vss.n264 268.425
R745 vss.n263 vss.n262 268.425
R746 vss.n972 vss.n130 268.425
R747 vss.n971 vss.n131 268.425
R748 vss.n954 vss.n953 268.425
R749 vss.n944 vss.n164 268.425
R750 vss.n277 vss.n230 268.425
R751 vss.n276 vss.n232 268.425
R752 vss.n778 vss.n721 268.425
R753 vss.n751 vss.n747 268.425
R754 vss.n762 vss.n761 268.425
R755 vss.n700 vss.n699 268.425
R756 vss.n705 vss.n704 268.425
R757 vss.n710 vss.n706 268.425
R758 vss.n665 vss.n663 268.274
R759 vss.n959 vss.n150 268.274
R760 vss.n252 vss.n249 268.274
R761 vss.n954 vss.n23 268.274
R762 vss.n944 vss.n943 268.274
R763 vss.n784 vss.n721 268.274
R764 vss.n700 vss.n653 268.274
R765 vss.n676 vss.n675 256.377
R766 vss.n674 vss.n673 256.377
R767 vss.n964 vss.n148 256.377
R768 vss.n147 vss.n146 256.377
R769 vss.n266 vss.n265 256.377
R770 vss.n264 vss.n263 256.377
R771 vss.n130 vss.n25 256.377
R772 vss.n972 vss.n971 256.377
R773 vss.n271 vss.n230 256.377
R774 vss.n277 vss.n276 256.377
R775 vss.n752 vss.n751 256.377
R776 vss.n761 vss.n747 256.377
R777 vss.n704 vss.n644 256.377
R778 vss.n706 vss.n705 256.377
R779 vss.n810 vss.n809 256
R780 vss.n216 vss.n215 256
R781 vss.n286 vss.n285 256
R782 vss.n951 vss.n161 256
R783 vss.n949 vss.n948 256
R784 vss.n777 vss.n728 256
R785 vss.n805 vss.n615 256
R786 vss.n115 vss.n40 251.859
R787 vss.n102 vss.n40 251.859
R788 vss.n86 vss.n85 251.859
R789 vss.n85 vss.n84 251.859
R790 vss.n69 vss.n61 251.859
R791 vss.n76 vss 251.859
R792 vss.n64 vss 251.859
R793 vss.n64 vss 251.859
R794 vss.n82 vss.n59 251.859
R795 vss.n71 vss.n59 251.859
R796 vss.n71 vss.n70 251.859
R797 vss.n70 vss.n69 251.859
R798 vss vss.n60 251.859
R799 vss.n77 vss 251.859
R800 vss.n77 vss 251.859
R801 vss vss.n76 251.859
R802 vss.n84 vss.n83 251.859
R803 vss.n83 vss.n82 251.859
R804 vss.n92 vss 251.859
R805 vss vss.n91 251.859
R806 vss.n91 vss 251.859
R807 vss.n60 vss 251.859
R808 vss.n104 vss.n98 251.859
R809 vss.n98 vss.n97 251.859
R810 vss.n97 vss.n54 251.859
R811 vss.n86 vss.n54 251.859
R812 vss vss.n53 251.859
R813 vss vss.n108 251.859
R814 vss.n108 vss 251.859
R815 vss.n92 vss 251.859
R816 vss.n103 vss.n102 251.859
R817 vss.n104 vss.n103 251.859
R818 vss vss.n41 251.859
R819 vss vss.n41 251.859
R820 vss.n53 vss 251.859
R821 vss.n116 vss.n115 251.859
R822 vss.n480 vss.n479 249.667
R823 vss.n922 vss.n295 216.847
R824 vss.n262 vss.n261 213.419
R825 vss.n145 vss.n144 213.407
R826 vss.n676 vss.n666 209.695
R827 vss.n641 vss.n637 209.695
R828 vss.n965 vss.n964 209.695
R829 vss.n267 vss.n266 209.695
R830 vss.n967 vss.n25 209.695
R831 vss.n202 vss.n131 209.695
R832 vss.n272 vss.n271 209.695
R833 vss.n236 vss.n232 209.695
R834 vss.n752 vss.n719 209.695
R835 vss.n762 vss.n738 209.695
R836 vss.n685 vss.n644 209.695
R837 vss.n711 vss.n710 209.695
R838 vss.n558 vss.n554 205.887
R839 vss.n518 vss.n299 188.065
R840 vss vss.n295 183.087
R841 vss.n925 vss.n924 151.014
R842 vss.n588 vss.n535 150.417
R843 vss.n484 vss.n328 150.417
R844 vss.n381 vss.n376 150.417
R845 vss.n465 vss.n464 150.417
R846 vss.n360 vss.n346 149.835
R847 vss.n360 vss 149.835
R848 vss.n348 vss.n346 149.835
R849 vss.n867 vss.n851 149.835
R850 vss.n852 vss.n851 149.835
R851 vss.n867 vss 149.835
R852 vss.n847 vss.n842 149.835
R853 vss.n871 vss.n842 149.835
R854 vss.n847 vss 149.835
R855 vss.n855 vss 149.835
R856 vss.n855 vss.n854 149.835
R857 vss.n862 vss.n854 149.835
R858 vss.n527 vss.n510 149.835
R859 vss.n527 vss 149.835
R860 vss.n511 vss.n510 149.835
R861 vss.n596 vss.n595 149.835
R862 vss.n595 vss 149.835
R863 vss.n597 vss.n596 149.835
R864 vss.n580 vss.n547 149.835
R865 vss.n560 vss.n552 149.835
R866 vss.n560 vss 149.835
R867 vss.n572 vss.n552 149.835
R868 vss.n556 vss.n553 149.835
R869 vss.n556 vss 149.835
R870 vss.n565 vss.n553 149.835
R871 vss.n520 vss.n514 149.835
R872 vss.n514 vss.n513 149.835
R873 vss.n513 vss 149.835
R874 vss.n591 vss 149.835
R875 vss.n591 vss.n502 149.835
R876 vss.n601 vss.n502 149.835
R877 vss.n830 vss.n818 149.835
R878 vss.n830 vss 149.835
R879 vss.n834 vss.n818 149.835
R880 vss.n828 vss.n825 149.835
R881 vss.n826 vss.n825 149.835
R882 vss.n828 vss 149.835
R883 vss.n857 vss.n309 149.835
R884 vss.n857 vss.n308 149.835
R885 vss vss.n308 149.835
R886 vss.n370 vss.n336 149.835
R887 vss.n370 vss 149.835
R888 vss.n337 vss.n336 149.835
R889 vss.n472 vss.n471 149.835
R890 vss.n434 vss.n407 149.835
R891 vss.n434 vss 149.835
R892 vss.n451 vss.n407 149.835
R893 vss.n421 vss.n417 149.835
R894 vss.n421 vss 149.835
R895 vss.n431 vss.n417 149.835
R896 vss.n355 vss.n351 149.835
R897 vss.n351 vss.n350 149.835
R898 vss.n350 vss 149.835
R899 vss.n366 vss.n339 149.835
R900 vss.n339 vss.n338 149.835
R901 vss.n338 vss 149.835
R902 vss.n440 vss.n439 149.835
R903 vss.n439 vss.n438 149.835
R904 vss.n438 vss 149.835
R905 vss.n476 vss.n385 149.835
R906 vss.n446 vss.n445 149.835
R907 vss.n419 vss 149.835
R908 vss.n426 vss.n419 149.835
R909 vss.n427 vss.n426 149.835
R910 vss.n359 vss.n348 149.459
R911 vss.n866 vss.n852 149.459
R912 vss.n872 vss.n871 149.459
R913 vss.n863 vss.n862 149.459
R914 vss.n526 vss.n511 149.459
R915 vss.n597 vss.n500 149.459
R916 vss.n572 vss.n571 149.459
R917 vss.n566 vss.n565 149.459
R918 vss.n521 vss.n520 149.459
R919 vss.n602 vss.n601 149.459
R920 vss.n835 vss.n834 149.459
R921 vss.n827 vss.n826 149.459
R922 vss.n874 vss.n309 149.459
R923 vss.n369 vss.n337 149.459
R924 vss.n452 vss.n451 149.459
R925 vss.n431 vss.n430 149.459
R926 vss.n356 vss.n355 149.459
R927 vss.n367 vss.n366 149.459
R928 vss.n440 vss.n406 149.459
R929 vss.n428 vss.n427 149.459
R930 vss.n119 vss.n118 138.59
R931 vss.n479 vss.n478 132.8
R932 vss.n465 vss 132.129
R933 vss.n588 vss 132.127
R934 vss vss.n328 132.127
R935 vss vss.n547 130.802
R936 vss.n472 vss 130.802
R937 vss.n446 vss 130.802
R938 vss.n478 vss.n477 120.001
R939 vss vss 118.966
R940 vss.n928 vss.n294 117.272
R941 vss.n601 vss.n600 117.001
R942 vss.n600 vss.n599 117.001
R943 vss.n592 vss.n591 117.001
R944 vss.n593 vss.n592 117.001
R945 vss.n520 vss.n519 117.001
R946 vss.n519 vss.n518 117.001
R947 vss.n513 vss.n506 117.001
R948 vss.n529 vss.n506 117.001
R949 vss.n565 vss.n564 117.001
R950 vss.n564 vss.n563 117.001
R951 vss.n557 vss.n556 117.001
R952 vss.n573 vss.n572 117.001
R953 vss.n574 vss.n573 117.001
R954 vss.n561 vss.n560 117.001
R955 vss.n562 vss.n561 117.001
R956 vss.n546 vss.n545 117.001
R957 vss.n545 vss.n540 117.001
R958 vss.n543 vss.n536 117.001
R959 vss.n543 vss.n541 117.001
R960 vss.n589 vss.n588 117.001
R961 vss.n590 vss.n589 117.001
R962 vss.n548 vss.n547 117.001
R963 vss.n575 vss.n548 117.001
R964 vss.n598 vss.n597 117.001
R965 vss.n599 vss.n598 117.001
R966 vss.n595 vss.n594 117.001
R967 vss.n594 vss.n593 117.001
R968 vss.n517 vss.n511 117.001
R969 vss.n518 vss.n517 117.001
R970 vss.n528 vss.n527 117.001
R971 vss.n529 vss.n528 117.001
R972 vss.n921 vss.n883 117.001
R973 vss.n888 vss.n883 117.001
R974 vss.n889 vss.n884 117.001
R975 vss.n916 vss.n889 117.001
R976 vss.n910 vss 117.001
R977 vss.n910 vss.n909 117.001
R978 vss.n903 vss.n902 117.001
R979 vss.n902 vss.n901 117.001
R980 vss vss.n896 117.001
R981 vss.n908 vss.n892 117.001
R982 vss.n909 vss.n908 117.001
R983 vss.n915 vss 117.001
R984 vss.n916 vss.n915 117.001
R985 vss vss.n882 117.001
R986 vss.n888 vss.n882 117.001
R987 vss.n297 vss.n294 117.001
R988 vss.n296 vss 117.001
R989 vss.n297 vss.n296 117.001
R990 vss.n754 vss.n753 117.001
R991 vss.n755 vss.n754 117.001
R992 vss.n749 vss.n748 117.001
R993 vss.n755 vss.n749 117.001
R994 vss.n780 vss.n779 117.001
R995 vss.n782 vss.n780 117.001
R996 vss.n784 vss.n783 117.001
R997 vss.n783 vss.n782 117.001
R998 vss.n679 vss.n678 117.001
R999 vss.n678 vss.n647 117.001
R1000 vss.n620 vss.n618 117.001
R1001 vss.n625 vss.n620 117.001
R1002 vss.n796 vss.n795 117.001
R1003 vss.n795 vss.n625 117.001
R1004 vss.n668 vss.n667 117.001
R1005 vss.n668 vss.n621 117.001
R1006 vss.n672 vss.n671 117.001
R1007 vss.n671 vss.n621 117.001
R1008 vss.n640 vss.n639 117.001
R1009 vss.n791 vss.n639 117.001
R1010 vss.n662 vss.n660 117.001
R1011 vss.n660 vss.n302 117.001
R1012 vss.n665 vss.n664 117.001
R1013 vss.n664 vss.n647 117.001
R1014 vss.n788 vss.n787 117.001
R1015 vss.n789 vss.n788 117.001
R1016 vss.n698 vss.n697 117.001
R1017 vss.n697 vss.n621 117.001
R1018 vss.n695 vss.n643 117.001
R1019 vss.n695 vss.n621 117.001
R1020 vss.n790 vss.n631 117.001
R1021 vss.n791 vss.n790 117.001
R1022 vss.n657 vss.n654 117.001
R1023 vss.n657 vss.n647 117.001
R1024 vss.n653 vss.n652 117.001
R1025 vss.n652 vss.n647 117.001
R1026 vss.n656 vss.n655 117.001
R1027 vss.n656 vss.n302 117.001
R1028 vss.n709 vss.n708 117.001
R1029 vss.n708 vss.n625 117.001
R1030 vss.n804 vss.n628 117.001
R1031 vss.n628 vss.n625 117.001
R1032 vss.n826 vss.n822 117.001
R1033 vss.n832 vss.n822 117.001
R1034 vss.n829 vss.n828 117.001
R1035 vss.n832 vss.n829 117.001
R1036 vss.n834 vss.n833 117.001
R1037 vss.n833 vss.n832 117.001
R1038 vss.n831 vss.n830 117.001
R1039 vss.n832 vss.n831 117.001
R1040 vss.n862 vss.n861 117.001
R1041 vss.n861 vss.n305 117.001
R1042 vss.n856 vss.n855 117.001
R1043 vss.n856 vss.n305 117.001
R1044 vss.n871 vss.n870 117.001
R1045 vss.n870 vss.n869 117.001
R1046 vss.n848 vss.n847 117.001
R1047 vss.n869 vss.n848 117.001
R1048 vss.n852 vss.n846 117.001
R1049 vss.n869 vss.n846 117.001
R1050 vss.n868 vss.n867 117.001
R1051 vss.n869 vss.n868 117.001
R1052 vss.n309 vss.n307 117.001
R1053 vss.n307 vss.n305 117.001
R1054 vss.n308 vss.n306 117.001
R1055 vss.n306 vss.n305 117.001
R1056 vss.n427 vss.n414 117.001
R1057 vss.n433 vss.n414 117.001
R1058 vss.n424 vss.n419 117.001
R1059 vss.n424 vss.n423 117.001
R1060 vss.n441 vss.n440 117.001
R1061 vss.n449 vss.n441 117.001
R1062 vss.n438 vss.n437 117.001
R1063 vss.n437 vss.n436 117.001
R1064 vss.n404 vss.n403 117.001
R1065 vss.n403 vss.n398 117.001
R1066 vss.n401 vss.n394 117.001
R1067 vss.n401 vss.n399 117.001
R1068 vss.n466 vss.n465 117.001
R1069 vss.n467 vss.n466 117.001
R1070 vss.n447 vss.n446 117.001
R1071 vss.n448 vss.n447 117.001
R1072 vss.n388 vss.n380 117.001
R1073 vss.n388 vss.n317 117.001
R1074 vss.n379 vss.n378 117.001
R1075 vss.n378 vss.n319 117.001
R1076 vss.n376 vss.n375 117.001
R1077 vss.n375 vss.n373 117.001
R1078 vss.n476 vss.n475 117.001
R1079 vss.n475 vss.n474 117.001
R1080 vss.n366 vss.n365 117.001
R1081 vss.n365 vss.n364 117.001
R1082 vss.n338 vss.n332 117.001
R1083 vss.n372 vss.n332 117.001
R1084 vss.n355 vss.n354 117.001
R1085 vss.n354 vss.n300 117.001
R1086 vss.n350 vss.n342 117.001
R1087 vss.n362 vss.n342 117.001
R1088 vss.n432 vss.n431 117.001
R1089 vss.n433 vss.n432 117.001
R1090 vss.n422 vss.n421 117.001
R1091 vss.n423 vss.n422 117.001
R1092 vss.n451 vss.n450 117.001
R1093 vss.n450 vss.n449 117.001
R1094 vss.n435 vss.n434 117.001
R1095 vss.n436 vss.n435 117.001
R1096 vss.n324 vss.n323 117.001
R1097 vss.n323 vss.n317 117.001
R1098 vss.n327 vss.n326 117.001
R1099 vss.n326 vss.n319 117.001
R1100 vss.n329 vss.n328 117.001
R1101 vss.n373 vss.n329 117.001
R1102 vss.n473 vss.n472 117.001
R1103 vss.n474 vss.n473 117.001
R1104 vss.n363 vss.n337 117.001
R1105 vss.n364 vss.n363 117.001
R1106 vss.n371 vss.n370 117.001
R1107 vss.n372 vss.n371 117.001
R1108 vss.n348 vss.n347 117.001
R1109 vss.n347 vss.n300 117.001
R1110 vss.n361 vss.n360 117.001
R1111 vss.n362 vss.n361 117.001
R1112 vss.n763 vss.n741 117.001
R1113 vss.n768 vss.n741 117.001
R1114 vss.n770 vss.n769 117.001
R1115 vss.n769 vss.n768 117.001
R1116 vss.n745 vss.n744 117.001
R1117 vss.n745 vss.n742 117.001
R1118 vss.n977 vss.n976 117.001
R1119 vss.n976 vss.n975 117.001
R1120 vss.n197 vss.n158 117.001
R1121 vss.n957 vss.n158 117.001
R1122 vss.n199 vss.n120 117.001
R1123 vss.n975 vss.n120 117.001
R1124 vss.n952 vss.n154 117.001
R1125 vss.n957 vss.n154 117.001
R1126 vss.n974 vss.n973 117.001
R1127 vss.n975 vss.n974 117.001
R1128 vss.n203 vss.n126 117.001
R1129 vss.n975 vss.n126 117.001
R1130 vss.n22 vss.n20 117.001
R1131 vss.n975 vss.n20 117.001
R1132 vss.n956 vss.n23 117.001
R1133 vss.n957 vss.n956 117.001
R1134 vss.n963 vss.n125 117.001
R1135 vss.n975 vss.n125 117.001
R1136 vss.n212 vss.n155 117.001
R1137 vss.n957 vss.n155 117.001
R1138 vss.n206 vss.n156 117.001
R1139 vss.n957 vss.n156 117.001
R1140 vss.n142 vss.n122 117.001
R1141 vss.n975 vss.n122 117.001
R1142 vss.n143 vss.n124 117.001
R1143 vss.n975 vss.n124 117.001
R1144 vss.n141 vss.n121 117.001
R1145 vss.n975 vss.n121 117.001
R1146 vss.n959 vss.n958 117.001
R1147 vss.n958 vss.n957 117.001
R1148 vss.n270 vss.n223 117.001
R1149 vss.n280 vss.n223 117.001
R1150 vss.n231 vss.n224 117.001
R1151 vss.n280 vss.n224 117.001
R1152 vss.n235 vss.n228 117.001
R1153 vss.n280 vss.n228 117.001
R1154 vss.n279 vss.n278 117.001
R1155 vss.n280 vss.n279 117.001
R1156 vss.n185 vss.n184 117.001
R1157 vss.n184 vss.n168 117.001
R1158 vss.n167 vss.n165 117.001
R1159 vss.n168 vss.n167 117.001
R1160 vss.n943 vss.n171 117.001
R1161 vss.n171 vss.n168 117.001
R1162 vss.n174 vss.n173 117.001
R1163 vss.n280 vss.n174 117.001
R1164 vss.n244 vss.n227 117.001
R1165 vss.n280 vss.n227 117.001
R1166 vss.n281 vss.n221 117.001
R1167 vss.n281 vss.n280 117.001
R1168 vss.n260 vss.n226 117.001
R1169 vss.n280 vss.n226 117.001
R1170 vss.n248 vss.n247 117.001
R1171 vss.n247 vss.n168 117.001
R1172 vss.n284 vss.n283 117.001
R1173 vss.n283 vss.n168 117.001
R1174 vss.n252 vss.n251 117.001
R1175 vss.n251 vss.n168 117.001
R1176 vss.n243 vss.n225 117.001
R1177 vss.n280 vss.n225 117.001
R1178 vss vss.n311 115.576
R1179 vss.n900 vss.n896 109.642
R1180 vss.n878 vss.n302 108.163
R1181 vss.n939 vss.n168 101.77
R1182 vss.n946 vss.n168 101.77
R1183 vss.n957 vss.n153 101.77
R1184 vss.n957 vss.n13 100.514
R1185 vss.n924 vss.n881 96.1003
R1186 vss.n781 vss.n716 90.9521
R1187 vss.n582 vss.n536 90.3534
R1188 vss.n587 vss.n536 90.3534
R1189 vss.n581 vss.n546 90.3534
R1190 vss.n576 vss.n546 90.3534
R1191 vss.n485 vss.n327 90.3534
R1192 vss.n327 vss.n314 90.3534
R1193 vss.n325 vss.n324 90.3534
R1194 vss.n324 vss.n313 90.3534
R1195 vss.n477 vss.n380 90.3534
R1196 vss.n384 vss.n380 90.3534
R1197 vss.n479 vss.n379 90.3534
R1198 vss.n382 vss.n379 90.3534
R1199 vss.n405 vss.n404 90.3534
R1200 vss.n404 vss.n395 90.3534
R1201 vss.n458 vss.n394 90.3534
R1202 vss.n463 vss.n394 90.3534
R1203 vss.n480 vss.n376 89.9911
R1204 vss.n969 vss.n123 89.6255
R1205 vss vss.n897 89.224
R1206 vss vss.n893 89.224
R1207 vss.n904 vss 89.224
R1208 vss.n904 vss.n903 89.224
R1209 vss vss.n885 89.224
R1210 vss vss.n914 89.224
R1211 vss.n914 vss.n892 89.224
R1212 vss.n897 vss.n892 89.224
R1213 vss.n885 vss 89.224
R1214 vss.n921 vss.n920 89.224
R1215 vss.n920 vss.n884 89.224
R1216 vss.n893 vss.n884 89.224
R1217 vss.n179 vss.n4 86.561
R1218 vss.n274 vss.n222 86.275
R1219 vss.n667 vss.n617 85.0829
R1220 vss.n667 vss.n635 85.0829
R1221 vss.n674 vss.n672 85.0829
R1222 vss.n796 vss.n637 85.0829
R1223 vss.n679 vss.n676 85.0829
R1224 vss.n147 vss.n142 85.0829
R1225 vss.n145 vss.n143 85.0829
R1226 vss.n964 vss.n963 85.0829
R1227 vss.n207 vss.n206 85.0829
R1228 vss.n206 vss.n9 85.0829
R1229 vss.n264 vss.n260 85.0829
R1230 vss.n259 vss.n248 85.0829
R1231 vss.n248 vss.n218 85.0829
R1232 vss.n266 vss.n244 85.0829
R1233 vss.n262 vss.n221 85.0829
R1234 vss.n199 vss.n131 85.0829
R1235 vss.n977 vss.n25 85.0829
R1236 vss.n953 vss.n952 85.0829
R1237 vss.n952 vss.n129 85.0829
R1238 vss.n973 vss.n972 85.0829
R1239 vss.n278 vss.n277 85.0829
R1240 vss.n186 vss.n185 85.0829
R1241 vss.n185 vss.n164 85.0829
R1242 vss.n271 vss.n270 85.0829
R1243 vss.n232 vss.n231 85.0829
R1244 vss.n748 vss.n747 85.0829
R1245 vss.n779 vss.n727 85.0829
R1246 vss.n779 vss.n778 85.0829
R1247 vss.n753 vss.n752 85.0829
R1248 vss.n763 vss.n762 85.0829
R1249 vss.n698 vss.n694 85.0829
R1250 vss.n699 vss.n698 85.0829
R1251 vss.n705 vss.n643 85.0829
R1252 vss.n654 vss.n644 85.0829
R1253 vss.n710 vss.n709 85.0829
R1254 vss.n683 vss.n662 84.9588
R1255 vss.n149 vss.n141 84.9588
R1256 vss.n253 vss.n243 84.9588
R1257 vss.n980 vss.n22 84.9588
R1258 vss.n941 vss.n173 84.9588
R1259 vss.n787 vss.n786 84.9588
R1260 vss.n689 vss.n655 84.9588
R1261 vss.n802 vss.n631 84.6953
R1262 vss.n640 vss.n632 84.6953
R1263 vss.n235 vss.n196 84.6953
R1264 vss.n204 vss.n203 84.6953
R1265 vss.n771 vss.n770 84.6953
R1266 vss.n939 vss.n179 83.5719
R1267 vss vss.n480 77.2563
R1268 vss.n975 vss.n119 71.1979
R1269 vss.n680 vss.n635 66.6518
R1270 vss.n961 vss.n9 66.6518
R1271 vss.n259 vss.n256 66.6518
R1272 vss.n129 vss.n24 66.6518
R1273 vss.n188 vss.n186 66.6518
R1274 vss.n733 vss.n727 66.6518
R1275 vss.n694 vss.n692 66.6518
R1276 vss.n798 vss.n797 64.7759
R1277 vss.n258 vss.n257 64.7759
R1278 vss.n984 vss.n10 64.7759
R1279 vss.n200 vss.n198 64.7759
R1280 vss.n937 vss.n187 64.7759
R1281 vss.n765 vss.n764 64.7759
R1282 vss.n693 vss.n629 64.7759
R1283 vss.n280 vss.n119 64.497
R1284 vss.n798 vss.n635 63.1207
R1285 vss.n259 vss.n258 63.1207
R1286 vss.n984 vss.n9 63.1207
R1287 vss.n198 vss.n129 63.1207
R1288 vss.n937 vss.n186 63.1207
R1289 vss.n765 vss.n727 63.1207
R1290 vss.n694 vss.n693 63.1207
R1291 vss.n877 vss.n303 61.4984
R1292 vss.n877 vss.n876 61.4984
R1293 vss.n681 vss.n680 61.2449
R1294 vss.n962 vss.n961 61.2449
R1295 vss.n256 vss.n255 61.2449
R1296 vss.n978 vss.n24 61.2449
R1297 vss.n188 vss.n172 61.2449
R1298 vss.n733 vss.n720 61.2449
R1299 vss.n692 vss.n691 61.2449
R1300 vss.n559 vss.n558 60.5013
R1301 vss.n581 vss.n580 59.4829
R1302 vss.n583 vss.n581 59.4829
R1303 vss.n583 vss.n582 59.4829
R1304 vss.n582 vss.n535 59.4829
R1305 vss.n471 vss.n325 59.4829
R1306 vss.n486 vss.n325 59.4829
R1307 vss.n486 vss.n485 59.4829
R1308 vss.n485 vss.n484 59.4829
R1309 vss.n385 vss.n384 59.4829
R1310 vss.n384 vss.n383 59.4829
R1311 vss.n383 vss.n382 59.4829
R1312 vss.n382 vss.n381 59.4829
R1313 vss.n445 vss.n395 59.4829
R1314 vss.n462 vss.n395 59.4829
R1315 vss.n463 vss.n462 59.4829
R1316 vss.n464 vss.n463 59.4829
R1317 vss.n797 vss.n796 58.5793
R1318 vss.n681 vss.n679 58.5793
R1319 vss.n143 vss.n10 58.5793
R1320 vss.n963 vss.n962 58.5793
R1321 vss.n255 vss.n244 58.5793
R1322 vss.n257 vss.n221 58.5793
R1323 vss.n200 vss.n199 58.5793
R1324 vss.n978 vss.n977 58.5793
R1325 vss.n270 vss.n172 58.5793
R1326 vss.n231 vss.n187 58.5793
R1327 vss.n753 vss.n720 58.5793
R1328 vss.n764 vss.n763 58.5793
R1329 vss.n691 vss.n654 58.5793
R1330 vss.n709 vss.n629 58.5793
R1331 vss.n672 vss.n635 54.2123
R1332 vss.n142 vss.n9 54.2123
R1333 vss.n260 vss.n259 54.2123
R1334 vss.n973 vss.n129 54.2123
R1335 vss.n278 vss.n186 54.2123
R1336 vss.n748 vss.n727 54.2123
R1337 vss.n694 vss.n643 54.2123
R1338 vss.n786 vss.n718 41.7862
R1339 vss.n724 vss.n718 41.7862
R1340 vss.n719 vss.n717 41.7862
R1341 vss.n756 vss.n717 41.7862
R1342 vss.n713 vss.n632 41.7862
R1343 vss.n792 vss.n713 41.7862
R1344 vss.n793 vss.n641 41.7862
R1345 vss.n793 vss.n792 41.7862
R1346 vss.n666 vss.n659 41.7862
R1347 vss.n687 vss.n659 41.7862
R1348 vss.n684 vss.n683 41.7862
R1349 vss.n687 vss.n684 41.7862
R1350 vss.n689 vss.n688 41.7862
R1351 vss.n688 vss.n687 41.7862
R1352 vss.n686 vss.n685 41.7862
R1353 vss.n687 vss.n686 41.7862
R1354 vss.n712 vss.n711 41.7862
R1355 vss.n792 vss.n712 41.7862
R1356 vss.n802 vss.n630 41.7862
R1357 vss.n792 vss.n630 41.7862
R1358 vss.n771 vss.n737 41.7862
R1359 vss.n767 vss.n737 41.7862
R1360 vss.n739 vss.n738 41.7862
R1361 vss.n740 vss.n739 41.7862
R1362 vss.n204 vss.n15 41.7862
R1363 vss.n982 vss.n15 41.7862
R1364 vss.n202 vss.n134 41.7862
R1365 vss.n969 vss.n134 41.7862
R1366 vss.n968 vss.n967 41.7862
R1367 vss.n969 vss.n968 41.7862
R1368 vss.n981 vss.n980 41.7862
R1369 vss.n982 vss.n981 41.7862
R1370 vss.n969 vss.n136 41.7862
R1371 vss.n966 vss.n965 41.7862
R1372 vss.n969 vss.n966 41.7862
R1373 vss.n149 vss.n18 41.7862
R1374 vss.n982 vss.n18 41.7862
R1375 vss.n196 vss.n177 41.7862
R1376 vss.n939 vss.n177 41.7862
R1377 vss.n941 vss.n940 41.7862
R1378 vss.n940 vss.n939 41.7862
R1379 vss.n273 vss.n272 41.7862
R1380 vss.n274 vss.n273 41.7862
R1381 vss.n237 vss.n236 41.7862
R1382 vss.n274 vss.n237 41.7862
R1383 vss.n253 vss.n181 41.7862
R1384 vss.n939 vss.n181 41.7862
R1385 vss.n268 vss.n267 41.7862
R1386 vss.n274 vss.n268 41.7862
R1387 vss.n274 vss.n239 41.7862
R1388 vss.n219 vss.n4 41.0949
R1389 vss vss.n576 40.4485
R1390 vss.n587 vss 40.4485
R1391 vss vss.n587 40.4485
R1392 vss vss.n313 40.4485
R1393 vss vss.n314 40.4485
R1394 vss vss.n314 40.4485
R1395 vss vss.n405 40.4485
R1396 vss vss.n458 40.4485
R1397 vss.n458 vss 40.4485
R1398 vss.n576 vss.n537 38.1445
R1399 vss.n490 vss.n313 38.1445
R1400 vss.n457 vss.n405 38.1445
R1401 vss.n144 vss.n136 37.7132
R1402 vss.n261 vss.n239 37.6975
R1403 vss.n927 vss.n926 34.4123
R1404 vss.n926 vss.n925 34.4123
R1405 vss.n714 vss.n293 34.4123
R1406 vss.n715 vss.n714 34.4123
R1407 vss.n733 vss.n732 34.4123
R1408 vss.n732 vss.n724 34.4123
R1409 vss.n723 vss.n721 34.4123
R1410 vss.n781 vss.n723 34.4123
R1411 vss.n757 vss.n751 34.4123
R1412 vss.n757 vss.n756 34.4123
R1413 vss.n680 vss.n650 34.4123
R1414 vss.n702 vss.n650 34.4123
R1415 vss.n798 vss.n624 34.4123
R1416 vss.n807 vss.n624 34.4123
R1417 vss.n673 vss.n626 34.4123
R1418 vss.n807 vss.n626 34.4123
R1419 vss.n675 vss.n651 34.4123
R1420 vss.n702 vss.n651 34.4123
R1421 vss.n663 vss.n649 34.4123
R1422 vss.n702 vss.n649 34.4123
R1423 vss.n809 vss.n808 34.4123
R1424 vss.n808 vss.n807 34.4123
R1425 vss.n806 vss.n805 34.4123
R1426 vss.n807 vss.n806 34.4123
R1427 vss.n701 vss.n700 34.4123
R1428 vss.n702 vss.n701 34.4123
R1429 vss.n692 vss.n648 34.4123
R1430 vss.n702 vss.n648 34.4123
R1431 vss.n693 vss.n623 34.4123
R1432 vss.n807 vss.n623 34.4123
R1433 vss.n704 vss.n703 34.4123
R1434 vss.n703 vss.n702 34.4123
R1435 vss.n706 vss.n622 34.4123
R1436 vss.n807 vss.n622 34.4123
R1437 vss.n766 vss.n765 34.4123
R1438 vss.n767 vss.n766 34.4123
R1439 vss.n743 vss.n728 34.4123
R1440 vss.n743 vss.n298 34.4123
R1441 vss.n761 vss.n760 34.4123
R1442 vss.n760 vss.n740 34.4123
R1443 vss.n24 vss.n14 34.4123
R1444 vss.n982 vss.n14 34.4123
R1445 vss.n198 vss.n19 34.4123
R1446 vss.n982 vss.n19 34.4123
R1447 vss.n971 vss.n970 34.4123
R1448 vss.n970 vss.n969 34.4123
R1449 vss.n133 vss.n130 34.4123
R1450 vss.n969 vss.n133 34.4123
R1451 vss.n955 vss.n954 34.4123
R1452 vss.n955 vss.n153 34.4123
R1453 vss.n161 vss.n160 34.4123
R1454 vss.n160 vss.n153 34.4123
R1455 vss.n961 vss.n16 34.4123
R1456 vss.n982 vss.n16 34.4123
R1457 vss.n984 vss.n983 34.4123
R1458 vss.n983 vss.n982 34.4123
R1459 vss.n146 vss.n139 34.4123
R1460 vss.n969 vss.n139 34.4123
R1461 vss.n148 vss.n135 34.4123
R1462 vss.n969 vss.n135 34.4123
R1463 vss.n151 vss.n150 34.4123
R1464 vss.n153 vss.n151 34.4123
R1465 vss.n215 vss.n214 34.4123
R1466 vss.n214 vss.n153 34.4123
R1467 vss.n188 vss.n176 34.4123
R1468 vss.n939 vss.n176 34.4123
R1469 vss.n938 vss.n937 34.4123
R1470 vss.n939 vss.n938 34.4123
R1471 vss.n948 vss.n947 34.4123
R1472 vss.n947 vss.n946 34.4123
R1473 vss.n945 vss.n944 34.4123
R1474 vss.n946 vss.n945 34.4123
R1475 vss.n234 vss.n230 34.4123
R1476 vss.n274 vss.n234 34.4123
R1477 vss.n276 vss.n275 34.4123
R1478 vss.n275 vss.n274 34.4123
R1479 vss.n256 vss.n178 34.4123
R1480 vss.n939 vss.n178 34.4123
R1481 vss.n258 vss.n180 34.4123
R1482 vss.n939 vss.n180 34.4123
R1483 vss.n285 vss.n169 34.4123
R1484 vss.n946 vss.n169 34.4123
R1485 vss.n249 vss.n170 34.4123
R1486 vss.n946 vss.n170 34.4123
R1487 vss.n265 vss.n238 34.4123
R1488 vss.n274 vss.n238 34.4123
R1489 vss.n263 vss.n241 34.4123
R1490 vss.n274 vss.n241 34.4123
R1491 vss.n61 vss.n31 32.5005
R1492 vss.n118 vss.n31 32.5005
R1493 vss vss.n48 32.5005
R1494 vss.n110 vss.n48 32.5005
R1495 vss vss.n47 32.5005
R1496 vss.n110 vss.n47 32.5005
R1497 vss.n70 vss.n33 32.5005
R1498 vss.n118 vss.n33 32.5005
R1499 vss vss.n46 32.5005
R1500 vss.n110 vss.n46 32.5005
R1501 vss.n83 vss.n34 32.5005
R1502 vss.n118 vss.n34 32.5005
R1503 vss.n59 vss.n30 32.5005
R1504 vss.n118 vss.n30 32.5005
R1505 vss vss.n49 32.5005
R1506 vss.n110 vss.n49 32.5005
R1507 vss.n85 vss.n29 32.5005
R1508 vss.n118 vss.n29 32.5005
R1509 vss vss.n50 32.5005
R1510 vss.n110 vss.n50 32.5005
R1511 vss vss.n45 32.5005
R1512 vss.n110 vss.n45 32.5005
R1513 vss.n54 vss.n35 32.5005
R1514 vss.n118 vss.n35 32.5005
R1515 vss vss.n44 32.5005
R1516 vss.n110 vss.n44 32.5005
R1517 vss.n103 vss.n36 32.5005
R1518 vss.n118 vss.n36 32.5005
R1519 vss.n98 vss.n28 32.5005
R1520 vss.n118 vss.n28 32.5005
R1521 vss.n109 vss 32.5005
R1522 vss.n110 vss.n109 32.5005
R1523 vss.n40 vss.n27 32.5005
R1524 vss.n118 vss.n27 32.5005
R1525 vss.n111 vss 32.5005
R1526 vss.n111 vss.n110 32.5005
R1527 vss vss.n42 32.5005
R1528 vss.n110 vss.n42 32.5005
R1529 vss.n117 vss.n116 32.5005
R1530 vss.n118 vss.n117 32.5005
R1531 vss.n939 vss.n119 25.5478
R1532 vss.n880 vss.n153 22.1973
R1533 vss.n63 vss.n62 19.5005
R1534 vss.n62 vss.n32 19.5005
R1535 vss.n68 vss.n67 19.5005
R1536 vss.n67 vss.n32 19.5005
R1537 vss.n75 vss.n74 19.5005
R1538 vss.n74 vss.n32 19.5005
R1539 vss.n81 vss.n80 19.5005
R1540 vss.n80 vss.n32 19.5005
R1541 vss.n58 vss.n57 19.5005
R1542 vss.n57 vss.n32 19.5005
R1543 vss.n90 vss.n89 19.5005
R1544 vss.n89 vss.n32 19.5005
R1545 vss.n96 vss.n95 19.5005
R1546 vss.n95 vss.n32 19.5005
R1547 vss.n107 vss.n106 19.5005
R1548 vss.n106 vss.n32 19.5005
R1549 vss.n101 vss.n100 19.5005
R1550 vss.n100 vss.n32 19.5005
R1551 vss.n114 vss.n113 19.5005
R1552 vss.n113 vss.n32 19.5005
R1553 vss.n39 vss.n37 19.5005
R1554 vss.n37 vss.n32 19.5005
R1555 vss.n946 vss.n119 18.8469
R1556 vss.n797 vss.n636 18.297
R1557 vss.n682 vss.n681 18.297
R1558 vss.n211 vss.n10 18.297
R1559 vss.n962 vss.n960 18.297
R1560 vss.n255 vss.n254 18.297
R1561 vss.n257 vss.n219 18.297
R1562 vss.n201 vss.n200 18.297
R1563 vss.n979 vss.n978 18.297
R1564 vss.n942 vss.n172 18.297
R1565 vss.n195 vss.n187 18.297
R1566 vss.n785 vss.n720 18.297
R1567 vss.n764 vss.n736 18.297
R1568 vss.n691 vss.n690 18.297
R1569 vss.n803 vss.n629 18.297
R1570 vss.n919 vss.n918 17.2064
R1571 vss.n918 vss.n917 17.2064
R1572 vss.n913 vss.n912 17.2064
R1573 vss.n912 vss.n890 17.2064
R1574 vss.n906 vss.n905 17.2064
R1575 vss.n906 vss.n895 17.2064
R1576 vss.n899 vss.n898 17.2064
R1577 vss.n923 vss.n922 17.2064
R1578 vss.n924 vss.n923 17.2064
R1579 vss.n280 vss.n222 15.4964
R1580 vss.n987 vss.n4 15.4704
R1581 vss.n119 vss.n17 12.9836
R1582 vss.n975 vss.n123 12.1459
R1583 vss.n683 vss.n682 8.08353
R1584 vss.n636 vss.n632 8.08353
R1585 vss.n960 vss.n149 8.08353
R1586 vss.n254 vss.n253 8.08353
R1587 vss.n980 vss.n979 8.08353
R1588 vss.n204 vss.n201 8.08353
R1589 vss.n942 vss.n941 8.08353
R1590 vss.n196 vss.n195 8.08353
R1591 vss.n786 vss.n785 8.08353
R1592 vss.n771 vss.n736 8.08353
R1593 vss.n690 vss.n689 8.08353
R1594 vss.n803 vss.n802 8.08353
R1595 vss.n839 vss.n838 6.69348
R1596 vss.n982 vss.n17 5.86382
R1597 vss.n901 vss.n900 5.84938
R1598 vss.n493 vss.n310 5.57706
R1599 vss.n499 vss 5.02361
R1600 vss.n312 vss 5.02361
R1601 vss.n312 vss 5.02361
R1602 vss.n455 vss 5.02361
R1603 vss.n568 vss 5.01717
R1604 vss.n569 vss 5.01717
R1605 vss.n501 vss 5.01717
R1606 vss.n501 vss 5.01717
R1607 vss.n524 vss 5.01717
R1608 vss.n524 vss 5.01717
R1609 vss.n837 vss 5.01717
R1610 vss.n817 vss 5.01717
R1611 vss.n853 vss 5.01717
R1612 vss.n853 vss 5.01717
R1613 vss.n864 vss 5.01717
R1614 vss.n864 vss 5.01717
R1615 vss.n418 vss 5.01717
R1616 vss.n418 vss 5.01717
R1617 vss.n454 vss 5.01717
R1618 vss.n454 vss 5.01717
R1619 vss.n349 vss 5.01717
R1620 vss.n349 vss 5.01717
R1621 vss.n357 vss 5.01717
R1622 vss.n357 vss 5.01717
R1623 vss.n567 vss.n495 4.99245
R1624 vss.n523 vss.n522 4.87797
R1625 vss.n512 vss.n498 4.50893
R1626 vss vss.n495 4.5005
R1627 vss.n608 vss.n496 4.5005
R1628 vss.n610 vss.n609 4.5005
R1629 vss.n605 vss.n604 4.5005
R1630 vss.n522 vss 4.5005
R1631 vss.n210 vss.n5 4.3205
R1632 vss.n985 vss.n8 3.27485
R1633 vss.n194 vss.n193 3.27485
R1634 vss.n936 vss.n189 3.27485
R1635 vss.n634 vss.n614 3.27485
R1636 vss.n799 vss.n613 3.27485
R1637 vss.n205 vss.n6 3.27485
R1638 vss.n735 vss.n734 3.27485
R1639 vss.n211 vss.n210 3.24353
R1640 vss.n636 vss.n618 3.08756
R1641 vss.n682 vss.n665 3.08756
R1642 vss.n212 vss.n211 3.08756
R1643 vss.n960 vss.n959 3.08756
R1644 vss.n254 vss.n252 3.08756
R1645 vss.n284 vss.n219 3.08756
R1646 vss.n201 vss.n197 3.08756
R1647 vss.n979 vss.n23 3.08756
R1648 vss.n943 vss.n942 3.08756
R1649 vss.n195 vss.n165 3.08756
R1650 vss.n785 vss.n784 3.08756
R1651 vss.n744 vss.n736 3.08756
R1652 vss.n690 vss.n653 3.08756
R1653 vss.n804 vss.n803 3.08756
R1654 vss.n289 vss 3.06629
R1655 vss.n191 vss 3.06629
R1656 vss.n813 vss 3.06629
R1657 vss.n478 vss 3.01226
R1658 vss.n0 vss 2.51601
R1659 vss.n841 vss.n840 2.46929
R1660 vss.n880 vss.n119 2.3703
R1661 vss.n43 vss.n39 2.35839
R1662 vss vss.n537 2.3045
R1663 vss.n490 vss 2.3045
R1664 vss vss.n457 2.3045
R1665 vss.n0 vss 2.11902
R1666 vss.n987 vss.n5 1.92736
R1667 vss.n616 vss 1.91991
R1668 vss.n217 vss 1.91991
R1669 vss.n163 vss 1.91991
R1670 vss.n525 vss.n521 1.8605
R1671 vss.n567 vss.n566 1.8605
R1672 vss.n571 vss.n570 1.8605
R1673 vss.n603 vss.n500 1.8605
R1674 vss.n526 vss.n525 1.8605
R1675 vss.n603 vss.n602 1.8605
R1676 vss.n836 vss.n835 1.8605
R1677 vss.n827 vss.n816 1.8605
R1678 vss.n874 vss.n873 1.8605
R1679 vss.n865 vss.n863 1.8605
R1680 vss.n873 vss.n872 1.8605
R1681 vss.n866 vss.n865 1.8605
R1682 vss.n453 vss.n406 1.8605
R1683 vss.n368 vss.n367 1.8605
R1684 vss.n358 vss.n356 1.8605
R1685 vss.n430 vss.n429 1.8605
R1686 vss.n453 vss.n452 1.8605
R1687 vss.n369 vss.n368 1.8605
R1688 vss.n359 vss.n358 1.8605
R1689 vss.n429 vss.n428 1.8605
R1690 vss.n494 vss.n493 1.79344
R1691 vss.n986 vss.n6 1.55665
R1692 vss.n986 vss.n985 1.55665
R1693 vss.n935 vss.n194 1.55665
R1694 vss.n936 vss.n935 1.55665
R1695 vss.n773 vss.n735 1.55665
R1696 vss.n800 vss.n634 1.55665
R1697 vss.n800 vss.n799 1.55665
R1698 vss.n290 vss.n205 1.43327
R1699 vss.n290 vss.n8 1.43327
R1700 vss.n193 vss.n192 1.43327
R1701 vss.n192 vss.n189 1.43327
R1702 vss.n734 vss.n292 1.43327
R1703 vss.n814 vss.n614 1.43327
R1704 vss.n814 vss.n613 1.43327
R1705 vss.n933 vss.n932 1.26772
R1706 vss.n982 vss.n13 1.25692
R1707 vss.n929 vss.n293 1.21955
R1708 vss.n840 vss.n839 1.14003
R1709 vss.n815 vss.n814 1.02854
R1710 vss.n606 vss.n605 0.99175
R1711 vss.n800 vss 0.946224
R1712 vss.n986 vss 0.946224
R1713 vss.n935 vss 0.946224
R1714 vss.n812 vss 0.905763
R1715 vss.n288 vss 0.905763
R1716 vss.n162 vss 0.905763
R1717 vss.n934 vss.n196 0.846996
R1718 vss.n934 vss.n204 0.846996
R1719 vss.n772 vss.n771 0.846996
R1720 vss.n802 vss.n801 0.846996
R1721 vss.n801 vss.n632 0.846996
R1722 vss vss 0.771099
R1723 vss.n537 vss.n497 0.715885
R1724 vss.n457 vss.n456 0.715885
R1725 vss.n491 vss.n311 0.715885
R1726 vss.n491 vss.n490 0.715885
R1727 vss.n775 vss 0.695143
R1728 vss.n258 vss.n6 0.664786
R1729 vss.n256 vss.n205 0.664786
R1730 vss.n985 vss.n984 0.664786
R1731 vss.n961 vss.n8 0.664786
R1732 vss.n198 vss.n194 0.664786
R1733 vss.n193 vss.n24 0.664786
R1734 vss.n937 vss.n936 0.664786
R1735 vss.n189 vss.n188 0.664786
R1736 vss.n765 vss.n735 0.664786
R1737 vss.n734 vss.n733 0.664786
R1738 vss.n931 vss 0.664786
R1739 vss.n693 vss.n634 0.664786
R1740 vss.n692 vss.n614 0.664786
R1741 vss.n799 vss.n798 0.664786
R1742 vss.n680 vss.n613 0.664786
R1743 vss.n731 vss 0.644695
R1744 vss vss 0.635531
R1745 vss.n927 vss.n295 0.582318
R1746 vss.n612 vss.n611 0.568833
R1747 vss.n989 vss.n3 0.52089
R1748 vss.n930 vss.n929 0.517167
R1749 vss vss 0.457722
R1750 vss.n633 vss 0.447211
R1751 vss.n7 vss 0.447211
R1752 vss.n190 vss 0.447211
R1753 vss.n192 vss 0.439349
R1754 vss.n290 vss 0.439349
R1755 vss.n814 vss 0.439349
R1756 vss.n606 vss.n496 0.418469
R1757 vss.n608 vss.n607 0.418469
R1758 vss.n611 vss.n610 0.414451
R1759 vss vss 0.406319
R1760 vss.n456 vss 0.405187
R1761 vss.n492 vss.n491 0.402844
R1762 vss.n607 vss.n497 0.401281
R1763 vss vss.n359 0.376971
R1764 vss vss.n866 0.376971
R1765 vss.n872 vss 0.376971
R1766 vss.n863 vss 0.376971
R1767 vss vss.n526 0.376971
R1768 vss vss.n500 0.376971
R1769 vss.n571 vss 0.376971
R1770 vss.n566 vss 0.376971
R1771 vss.n521 vss 0.376971
R1772 vss.n602 vss 0.376971
R1773 vss.n835 vss 0.376971
R1774 vss.n810 vss.n617 0.376971
R1775 vss.n216 vss.n207 0.376971
R1776 vss.n286 vss.n218 0.376971
R1777 vss.n953 vss.n951 0.376971
R1778 vss.n949 vss.n164 0.376971
R1779 vss.n778 vss.n777 0.376971
R1780 vss.n699 vss.n615 0.376971
R1781 vss vss.n827 0.376971
R1782 vss vss.n874 0.376971
R1783 vss vss.n369 0.376971
R1784 vss.n452 vss 0.376971
R1785 vss.n430 vss 0.376971
R1786 vss.n356 vss 0.376971
R1787 vss.n367 vss 0.376971
R1788 vss vss.n406 0.376971
R1789 vss.n478 vss.n311 0.376971
R1790 vss.n428 vss 0.376971
R1791 vss.n499 vss.n497 0.376281
R1792 vss.n456 vss.n455 0.376281
R1793 vss.n491 vss.n312 0.376281
R1794 vss.n990 vss.n2 0.367058
R1795 vss.n605 vss.n498 0.35393
R1796 vss.n773 vss 0.342762
R1797 vss.n633 vss.n616 0.321553
R1798 vss.n813 vss.n812 0.321553
R1799 vss.n217 vss.n7 0.321553
R1800 vss.n289 vss.n288 0.321553
R1801 vss.n190 vss.n163 0.321553
R1802 vss.n191 vss.n162 0.321553
R1803 vss.n774 vss 0.318384
R1804 vss.n43 vss.n2 0.304262
R1805 vss.n610 vss.n496 0.301281
R1806 vss.n609 vss.n608 0.301281
R1807 vss.n612 vss.n494 0.250766
R1808 vss.n840 vss.n612 0.250595
R1809 vss.n775 vss.n774 0.228964
R1810 vss.n839 vss.n815 0.226195
R1811 vss.n2 vss.n1 0.218382
R1812 vss vss.n836 0.208833
R1813 vss.n1 vss.n0 0.188289
R1814 vss.n812 vss.n811 0.186355
R1815 vss.n288 vss.n287 0.186355
R1816 vss.n950 vss.n162 0.186355
R1817 vss.n989 vss.n988 0.181262
R1818 vss.n800 vss.n633 0.171553
R1819 vss.n986 vss.n7 0.171553
R1820 vss.n935 vss.n190 0.171553
R1821 vss.n291 vss 0.166889
R1822 vss vss.n603 0.166125
R1823 vss.n368 vss 0.166125
R1824 vss.n570 vss 0.164562
R1825 vss.n525 vss 0.164562
R1826 vss.n865 vss 0.164562
R1827 vss.n453 vss 0.164562
R1828 vss.n358 vss 0.164562
R1829 vss.n811 vss.n616 0.158395
R1830 vss.n287 vss.n217 0.158395
R1831 vss.n950 vss.n163 0.158395
R1832 vss.n816 vss.n815 0.14931
R1833 vss.n290 vss.n289 0.145237
R1834 vss.n192 vss.n191 0.145237
R1835 vss.n814 vss.n813 0.145237
R1836 vss.n836 vss.n817 0.139389
R1837 vss.n990 vss 0.138431
R1838 vss.n811 vss.n810 0.133357
R1839 vss.n287 vss.n216 0.133357
R1840 vss.n287 vss.n286 0.133357
R1841 vss.n951 vss.n950 0.133357
R1842 vss.n950 vss.n949 0.133357
R1843 vss.n777 vss.n776 0.133357
R1844 vss.n811 vss.n615 0.133357
R1845 vss.n731 vss 0.126904
R1846 vss vss.n933 0.124938
R1847 vss vss.n291 0.123766
R1848 vss.n1 vss 0.111032
R1849 vss.n838 vss.n816 0.110619
R1850 vss.n568 vss.n567 0.109875
R1851 vss.n570 vss.n569 0.109875
R1852 vss.n603 vss.n501 0.109875
R1853 vss.n525 vss.n524 0.109875
R1854 vss.n865 vss.n864 0.109875
R1855 vss.n429 vss.n418 0.109875
R1856 vss.n454 vss.n453 0.109875
R1857 vss.n358 vss.n357 0.109875
R1858 vss.n609 vss 0.109094
R1859 vss.n729 vss 0.10256
R1860 vss.n368 vss.n310 0.0903438
R1861 vss.n853 vss.n841 0.0860255
R1862 vss.n773 vss.n772 0.0803611
R1863 vss.n607 vss.n606 0.0780862
R1864 vss.n493 vss.n492 0.0780862
R1865 vss vss 0.0768081
R1866 vss.n292 vss 0.0759438
R1867 vss.n837 vss 0.0699444
R1868 vss.n817 vss 0.0699444
R1869 vss.n776 vss.n731 0.0677619
R1870 vss.n815 vss 0.065907
R1871 vss.n987 vss.n986 0.0651358
R1872 vss.n935 vss.n934 0.0651358
R1873 vss.n934 vss 0.0651358
R1874 vss.n801 vss.n800 0.0651358
R1875 vss.n801 vss 0.0651358
R1876 vss.n774 vss.n773 0.0624048
R1877 vss.n3 vss 0.0620278
R1878 vss.n776 vss.n775 0.0576429
R1879 vss.n988 vss 0.0572671
R1880 vss vss.n568 0.0551875
R1881 vss.n569 vss 0.0551875
R1882 vss vss.n853 0.0551875
R1883 vss.n864 vss 0.0551875
R1884 vss.n418 vss 0.0551875
R1885 vss vss.n454 0.0551875
R1886 vss vss.n349 0.0551875
R1887 vss.n357 vss 0.0551875
R1888 vss vss.n730 0.0524663
R1889 vss.n455 vss 0.0434688
R1890 vss vss.n312 0.0434688
R1891 vss.n730 vss 0.0433241
R1892 vss.n933 vss.n290 0.042429
R1893 vss.n730 vss.n729 0.0417809
R1894 vss.n729 vss.n292 0.0416985
R1895 vss.n604 vss.n499 0.0395625
R1896 vss.n522 vss.n498 0.0354764
R1897 vss.n611 vss.n495 0.034875
R1898 vss vss.n990 0.0326121
R1899 vss.n932 vss.n931 0.0316884
R1900 vss.n524 vss.n523 0.0309688
R1901 vss vss.n512 0.0301875
R1902 vss.n932 vss.n291 0.0294694
R1903 vss.n838 vss.n837 0.0292698
R1904 vss.n512 vss.n501 0.0255
R1905 vss.n523 vss 0.0247187
R1906 vss.n873 vss.n841 0.0233551
R1907 vss.n349 vss.n310 0.0200312
R1908 vss.n772 vss.n3 0.0188333
R1909 vss.n930 vss.n292 0.0120878
R1910 vss vss.n989 0.00952437
R1911 vss.n988 vss.n987 0.00836871
R1912 vss.n494 vss 0.00513139
R1913 vss.n604 vss 0.00440625
R1914 vss.n492 vss 0.00284375
R1915 vss.n931 vss.n930 0.000993097
R1916 vdd.n600 vdd.n580 5809.41
R1917 vdd.n643 vdd.n600 5809.41
R1918 vdd.n682 vdd.n501 5809.41
R1919 vdd.n501 vdd.n498 5809.41
R1920 vdd.n726 vdd.n691 5809.41
R1921 vdd.n726 vdd.n692 5809.41
R1922 vdd.n729 vdd.n728 5809.41
R1923 vdd.n728 vdd.n483 5809.41
R1924 vdd.n497 vdd.n495 5809.41
R1925 vdd.n684 vdd.n495 5809.41
R1926 vdd.n787 vdd.n39 5809.41
R1927 vdd.n787 vdd.n40 5809.41
R1928 vdd.n815 vdd.n16 5809.41
R1929 vdd.n16 vdd.n13 5809.41
R1930 vdd.n627 vdd.n624 5784.71
R1931 vdd.n628 vdd.n627 5784.71
R1932 vdd.n553 vdd.n487 5784.71
R1933 vdd.n551 vdd.n487 5784.71
R1934 vdd.n713 vdd.n708 5784.71
R1935 vdd.n709 vdd.n708 5784.71
R1936 vdd.n706 vdd.n697 5784.71
R1937 vdd.n706 vdd.n698 5784.71
R1938 vdd.n689 vdd.n489 5784.71
R1939 vdd.n689 vdd.n490 5784.71
R1940 vdd.n70 vdd.n55 5784.71
R1941 vdd.n57 vdd.n55 5784.71
R1942 vdd.n807 vdd.n26 5784.71
R1943 vdd.n809 vdd.n26 5784.71
R1944 vdd.n597 vdd.n585 4912.94
R1945 vdd.n589 vdd.n585 4912.94
R1946 vdd.n597 vdd.n586 4912.94
R1947 vdd.n640 vdd.n603 4912.94
R1948 vdd.n640 vdd.n639 4912.94
R1949 vdd.n639 vdd.n604 4912.94
R1950 vdd.n604 vdd.n603 4912.94
R1951 vdd.n674 vdd.n513 4912.94
R1952 vdd.n674 vdd.n514 4912.94
R1953 vdd.n513 vdd.n509 4912.94
R1954 vdd.n514 vdd.n509 4912.94
R1955 vdd.n506 vdd.n505 4912.94
R1956 vdd.n677 vdd.n505 4912.94
R1957 vdd.n676 vdd.n506 4912.94
R1958 vdd.n677 vdd.n676 4912.94
R1959 vdd.n743 vdd.n469 4912.94
R1960 vdd.n722 vdd.n469 4912.94
R1961 vdd.n743 vdd.n470 4912.94
R1962 vdd.n722 vdd.n470 4912.94
R1963 vdd.n741 vdd.n472 4912.94
R1964 vdd.n720 vdd.n472 4912.94
R1965 vdd.n741 vdd.n473 4912.94
R1966 vdd.n720 vdd.n473 4912.94
R1967 vdd.n796 vdd.n792 4912.94
R1968 vdd.n794 vdd.n792 4912.94
R1969 vdd.n53 vdd.n52 4912.94
R1970 vdd.n76 vdd.n52 4912.94
R1971 vdd.n73 vdd.n53 4912.94
R1972 vdd.n76 vdd.n73 4912.94
R1973 vdd.n794 vdd.n793 4849.41
R1974 vdd.n613 vdd.n612 4207.06
R1975 vdd.n579 vdd.n577 4207.06
R1976 vdd.n646 vdd.n577 4207.06
R1977 vdd.n636 vdd.n613 4207.06
R1978 vdd.n561 vdd.n541 4207.06
R1979 vdd.n541 vdd.n540 4207.06
R1980 vdd.n665 vdd.n536 4207.06
R1981 vdd.n665 vdd.n664 4207.06
R1982 vdd.n747 vdd.n460 4207.06
R1983 vdd.n749 vdd.n460 4207.06
R1984 vdd.n755 vdd.n456 4207.06
R1985 vdd.n456 vdd.n452 4207.06
R1986 vdd.n522 vdd.n519 4207.06
R1987 vdd.n523 vdd.n522 4207.06
R1988 vdd.n667 vdd.n524 4207.06
R1989 vdd.n668 vdd.n667 4207.06
R1990 vdd.n475 vdd.n465 4207.06
R1991 vdd.n475 vdd.n463 4207.06
R1992 vdd.n757 vdd.n450 4207.06
R1993 vdd.n453 vdd.n450 4207.06
R1994 vdd.n791 vdd.n33 4207.06
R1995 vdd.n803 vdd.n791 4207.06
R1996 vdd.n67 vdd.n61 4207.06
R1997 vdd.n61 vdd.n59 4207.06
R1998 vdd.n775 vdd.n80 4207.06
R1999 vdd.n776 vdd.n775 4207.06
R2000 vdd.n624 vdd.n616 4020
R2001 vdd.n628 vdd.n582 4020
R2002 vdd.n553 vdd.n500 4020
R2003 vdd.n551 vdd.n550 4020
R2004 vdd.n713 vdd.n712 4020
R2005 vdd.n710 vdd.n709 4020
R2006 vdd.n697 vdd.n482 4020
R2007 vdd.n700 vdd.n698 4020
R2008 vdd.n510 vdd.n489 4020
R2009 vdd.n494 vdd.n490 4020
R2010 vdd.n70 vdd.n44 4020
R2011 vdd.n57 vdd.n45 4020
R2012 vdd.n807 vdd.n15 4020
R2013 vdd.n810 vdd.n809 4020
R2014 vdd.n616 vdd.n580 3998.82
R2015 vdd.n643 vdd.n582 3998.82
R2016 vdd.n682 vdd.n500 3998.82
R2017 vdd.n550 vdd.n498 3998.82
R2018 vdd.n712 vdd.n691 3998.82
R2019 vdd.n710 vdd.n692 3998.82
R2020 vdd.n729 vdd.n482 3998.82
R2021 vdd.n700 vdd.n483 3998.82
R2022 vdd.n510 vdd.n497 3998.82
R2023 vdd.n684 vdd.n494 3998.82
R2024 vdd.n44 vdd.n39 3998.82
R2025 vdd.n45 vdd.n40 3998.82
R2026 vdd.n815 vdd.n15 3998.82
R2027 vdd.n810 vdd.n13 3998.82
R2028 vdd.n818 vdd.n10 3734.12
R2029 vdd.n612 vdd.n611 3409.41
R2030 vdd.n611 vdd.n579 3409.41
R2031 vdd.n636 vdd.n576 3409.41
R2032 vdd.n646 vdd.n576 3409.41
R2033 vdd.n562 vdd.n561 3409.41
R2034 vdd.n562 vdd.n536 3409.41
R2035 vdd.n540 vdd.n537 3409.41
R2036 vdd.n664 vdd.n537 3409.41
R2037 vdd.n747 vdd.n455 3409.41
R2038 vdd.n755 vdd.n455 3409.41
R2039 vdd.n750 vdd.n749 3409.41
R2040 vdd.n750 vdd.n452 3409.41
R2041 vdd.n519 vdd.n518 3409.41
R2042 vdd.n524 vdd.n518 3409.41
R2043 vdd.n669 vdd.n523 3409.41
R2044 vdd.n669 vdd.n668 3409.41
R2045 vdd.n465 vdd.n449 3409.41
R2046 vdd.n757 vdd.n449 3409.41
R2047 vdd.n733 vdd.n463 3409.41
R2048 vdd.n733 vdd.n453 3409.41
R2049 vdd.n33 vdd.n9 3409.41
R2050 vdd.n818 vdd.n9 3409.41
R2051 vdd.n803 vdd.n802 3409.41
R2052 vdd.n802 vdd.n12 3409.41
R2053 vdd.n67 vdd.n48 3409.41
R2054 vdd.n80 vdd.n48 3409.41
R2055 vdd.n59 vdd.n49 3409.41
R2056 vdd.n776 vdd.n49 3409.41
R2057 vdd.n618 vdd.n616 1789.41
R2058 vdd.n618 vdd.n582 1789.41
R2059 vdd.n433 vdd.n407 1789.41
R2060 vdd.n407 vdd.n403 1789.41
R2061 vdd.n433 vdd.n408 1789.41
R2062 vdd.n408 vdd.n403 1789.41
R2063 vdd.n406 vdd.n400 1789.41
R2064 vdd.n435 vdd.n400 1789.41
R2065 vdd.n406 vdd.n401 1789.41
R2066 vdd.n435 vdd.n401 1789.41
R2067 vdd.n416 vdd.n411 1789.41
R2068 vdd.n425 vdd.n411 1789.41
R2069 vdd.n416 vdd.n412 1789.41
R2070 vdd.n425 vdd.n412 1789.41
R2071 vdd.n418 vdd.n414 1789.41
R2072 vdd.n423 vdd.n418 1789.41
R2073 vdd.n419 vdd.n414 1789.41
R2074 vdd.n423 vdd.n419 1789.41
R2075 vdd.n153 vdd.n141 1789.41
R2076 vdd.n150 vdd.n141 1789.41
R2077 vdd.n153 vdd.n142 1789.41
R2078 vdd.n159 vdd.n136 1789.41
R2079 vdd.n156 vdd.n136 1789.41
R2080 vdd.n159 vdd.n137 1789.41
R2081 vdd.n156 vdd.n137 1789.41
R2082 vdd.n123 vdd.n94 1789.41
R2083 vdd.n123 vdd.n95 1789.41
R2084 vdd.n163 vdd.n87 1789.41
R2085 vdd.n134 vdd.n87 1789.41
R2086 vdd.n116 vdd.n97 1789.41
R2087 vdd.n119 vdd.n97 1789.41
R2088 vdd.n116 vdd.n98 1789.41
R2089 vdd.n119 vdd.n98 1789.41
R2090 vdd.n113 vdd.n102 1789.41
R2091 vdd.n110 vdd.n103 1789.41
R2092 vdd.n113 vdd.n103 1789.41
R2093 vdd.n549 vdd.n500 1789.41
R2094 vdd.n550 vdd.n549 1789.41
R2095 vdd.n712 vdd.n711 1789.41
R2096 vdd.n711 vdd.n710 1789.41
R2097 vdd.n701 vdd.n482 1789.41
R2098 vdd.n701 vdd.n700 1789.41
R2099 vdd.n511 vdd.n510 1789.41
R2100 vdd.n511 vdd.n494 1789.41
R2101 vdd.n782 vdd.n44 1789.41
R2102 vdd.n782 vdd.n45 1789.41
R2103 vdd.n811 vdd.n15 1789.41
R2104 vdd.n811 vdd.n810 1789.41
R2105 vdd.n203 vdd.n188 1789.41
R2106 vdd.n210 vdd.n188 1789.41
R2107 vdd.n203 vdd.n189 1789.41
R2108 vdd.n210 vdd.n189 1789.41
R2109 vdd.n219 vdd.n181 1789.41
R2110 vdd.n200 vdd.n181 1789.41
R2111 vdd.n219 vdd.n182 1789.41
R2112 vdd.n200 vdd.n182 1789.41
R2113 vdd.n331 vdd.n324 1789.41
R2114 vdd.n324 vdd.n322 1789.41
R2115 vdd.n343 vdd.n176 1789.41
R2116 vdd.n345 vdd.n176 1789.41
R2117 vdd.n305 vdd.n286 1789.41
R2118 vdd.n305 vdd.n287 1789.41
R2119 vdd.n319 vdd.n245 1789.41
R2120 vdd.n319 vdd.n246 1789.41
R2121 vdd.n279 vdd.n251 1789.41
R2122 vdd.n308 vdd.n251 1789.41
R2123 vdd.n279 vdd.n252 1789.41
R2124 vdd.n308 vdd.n252 1789.41
R2125 vdd.n271 vdd.n263 1789.41
R2126 vdd.n263 vdd.n258 1789.41
R2127 vdd.n271 vdd.n264 1789.41
R2128 vdd.n264 vdd.n258 1789.41
R2129 vdd.n205 vdd.n191 1789.41
R2130 vdd.n208 vdd.n191 1789.41
R2131 vdd.n205 vdd.n192 1789.41
R2132 vdd.n208 vdd.n192 1789.41
R2133 vdd.n194 vdd.n179 1789.41
R2134 vdd.n199 vdd.n194 1789.41
R2135 vdd.n195 vdd.n179 1789.41
R2136 vdd.n199 vdd.n195 1789.41
R2137 vdd.n323 vdd.n242 1789.41
R2138 vdd.n333 vdd.n242 1789.41
R2139 vdd.n238 vdd.n222 1789.41
R2140 vdd.n238 vdd.n178 1789.41
R2141 vdd.n281 vdd.n254 1789.41
R2142 vdd.n284 vdd.n254 1789.41
R2143 vdd.n281 vdd.n255 1789.41
R2144 vdd.n284 vdd.n255 1789.41
R2145 vdd.n273 vdd.n259 1789.41
R2146 vdd.n276 vdd.n259 1789.41
R2147 vdd.n273 vdd.n260 1789.41
R2148 vdd.n276 vdd.n260 1789.41
R2149 vdd.n389 vdd.n363 1789.41
R2150 vdd.n363 vdd.n359 1789.41
R2151 vdd.n389 vdd.n364 1789.41
R2152 vdd.n364 vdd.n359 1789.41
R2153 vdd.n362 vdd.n356 1789.41
R2154 vdd.n391 vdd.n356 1789.41
R2155 vdd.n362 vdd.n357 1789.41
R2156 vdd.n391 vdd.n357 1789.41
R2157 vdd.n372 vdd.n367 1789.41
R2158 vdd.n381 vdd.n367 1789.41
R2159 vdd.n372 vdd.n368 1789.41
R2160 vdd.n381 vdd.n368 1789.41
R2161 vdd.n374 vdd.n370 1789.41
R2162 vdd.n379 vdd.n374 1789.41
R2163 vdd.n375 vdd.n370 1789.41
R2164 vdd.n379 vdd.n375 1789.41
R2165 vdd.n598 vdd.n584 1534.21
R2166 vdd.n122 vdd.n120 1315.04
R2167 vdd.n89 vdd.n86 1231.76
R2168 vdd.n90 vdd.n89 1231.76
R2169 vdd.n129 vdd.n128 1231.76
R2170 vdd.n128 vdd.n92 1231.76
R2171 vdd.n224 vdd.n223 1231.76
R2172 vdd.n223 vdd.n175 1231.76
R2173 vdd.n326 vdd.n226 1231.76
R2174 vdd.n326 vdd.n325 1231.76
R2175 vdd.n295 vdd.n294 1231.76
R2176 vdd.n294 vdd.n293 1231.76
R2177 vdd.n300 vdd.n289 1231.76
R2178 vdd.n300 vdd.n290 1231.76
R2179 vdd.n234 vdd.n231 1231.76
R2180 vdd.n234 vdd.n233 1231.76
R2181 vdd.n335 vdd.n230 1231.76
R2182 vdd.n335 vdd.n334 1231.76
R2183 vdd.n589 vdd.n588 1189.42
R2184 vdd.n611 vdd.n610 797.648
R2185 vdd.n610 vdd.n576 797.648
R2186 vdd.n563 vdd.n562 797.648
R2187 vdd.n563 vdd.n537 797.648
R2188 vdd.n751 vdd.n455 797.648
R2189 vdd.n751 vdd.n750 797.648
R2190 vdd.n670 vdd.n518 797.648
R2191 vdd.n670 vdd.n669 797.648
R2192 vdd.n734 vdd.n449 797.648
R2193 vdd.n734 vdd.n733 797.648
R2194 vdd.n801 vdd.n9 797.648
R2195 vdd.n802 vdd.n801 797.648
R2196 vdd.n780 vdd.n48 797.648
R2197 vdd.n780 vdd.n49 797.648
R2198 vdd.n129 vdd.n94 557.648
R2199 vdd.n130 vdd.n129 557.648
R2200 vdd.n130 vdd.n86 557.648
R2201 vdd.n163 vdd.n86 557.648
R2202 vdd.n95 vdd.n92 557.648
R2203 vdd.n132 vdd.n92 557.648
R2204 vdd.n132 vdd.n90 557.648
R2205 vdd.n134 vdd.n90 557.648
R2206 vdd.n331 vdd.n226 557.648
R2207 vdd.n341 vdd.n226 557.648
R2208 vdd.n341 vdd.n224 557.648
R2209 vdd.n343 vdd.n224 557.648
R2210 vdd.n325 vdd.n322 557.648
R2211 vdd.n325 vdd.n228 557.648
R2212 vdd.n228 vdd.n175 557.648
R2213 vdd.n345 vdd.n175 557.648
R2214 vdd.n289 vdd.n286 557.648
R2215 vdd.n297 vdd.n289 557.648
R2216 vdd.n297 vdd.n295 557.648
R2217 vdd.n295 vdd.n245 557.648
R2218 vdd.n290 vdd.n287 557.648
R2219 vdd.n291 vdd.n290 557.648
R2220 vdd.n293 vdd.n291 557.648
R2221 vdd.n293 vdd.n246 557.648
R2222 vdd.n323 vdd.n230 557.648
R2223 vdd.n339 vdd.n230 557.648
R2224 vdd.n339 vdd.n231 557.648
R2225 vdd.n231 vdd.n222 557.648
R2226 vdd.n334 vdd.n333 557.648
R2227 vdd.n334 vdd.n229 557.648
R2228 vdd.n233 vdd.n229 557.648
R2229 vdd.n233 vdd.n178 557.648
R2230 vdd vdd.n587 524.352
R2231 vdd.n596 vdd.n587 524.068
R2232 vdd.n5 vdd.n4 486.526
R2233 vdd.n590 vdd 478.745
R2234 vdd.n599 vdd.n598 473.772
R2235 vdd.n596 vdd.n595 473.219
R2236 vdd.n621 vdd.n620 447.06
R2237 vdd.n681 vdd.n680 447.06
R2238 vdd.n725 vdd.n716 447.06
R2239 vdd.n699 vdd.n485 447.06
R2240 vdd.n685 vdd.n493 447.06
R2241 vdd.n786 vdd.n785 447.06
R2242 vdd.n24 vdd.n23 447.06
R2243 vdd.n623 vdd.n614 444.515
R2244 vdd.n555 vdd.n554 444.515
R2245 vdd.n714 vdd.n696 444.515
R2246 vdd.n705 vdd.n704 444.515
R2247 vdd.n688 vdd.n687 444.515
R2248 vdd.n62 vdd.n42 444.515
R2249 vdd.n35 vdd.n27 444.515
R2250 vdd.n623 vdd.n622 428.8
R2251 vdd.n554 vdd.n502 428.8
R2252 vdd.n715 vdd.n714 428.8
R2253 vdd.n704 vdd.n703 428.8
R2254 vdd.n687 vdd.n686 428.8
R2255 vdd.n784 vdd.n42 428.8
R2256 vdd.n27 vdd.n25 428.8
R2257 vdd.n622 vdd.n621 426.541
R2258 vdd.n681 vdd.n502 426.541
R2259 vdd.n716 vdd.n715 426.541
R2260 vdd.n703 vdd.n699 426.541
R2261 vdd.n686 vdd.n685 426.541
R2262 vdd.n785 vdd.n784 426.541
R2263 vdd.n25 vdd.n24 426.541
R2264 vdd.n819 vdd.n8 378.38
R2265 vdd.n635 vdd.n574 363.671
R2266 vdd.n565 vdd.n538 363.671
R2267 vdd.n461 vdd.n459 363.671
R2268 vdd.n474 vdd.n447 363.671
R2269 vdd.n520 vdd.n517 363.671
R2270 vdd.n66 vdd.n50 363.671
R2271 vdd.n34 vdd.n7 363.671
R2272 vdd.n648 vdd.n647 363.295
R2273 vdd.n663 vdd.n662 363.295
R2274 vdd.n717 vdd.n444 363.295
R2275 vdd.n759 vdd.n758 363.295
R2276 vdd.n568 vdd.n567 363.295
R2277 vdd.n773 vdd.n772 363.295
R2278 vdd.n820 vdd.n819 363.295
R2279 vdd.n635 vdd.n634 362.37
R2280 vdd.n556 vdd.n538 362.37
R2281 vdd.n521 vdd.n520 362.37
R2282 vdd.n467 vdd.n461 362.37
R2283 vdd.n476 vdd.n474 362.37
R2284 vdd.n37 vdd.n34 362.37
R2285 vdd.n66 vdd.n65 362.37
R2286 vdd.n647 vdd.n575 361.584
R2287 vdd.n663 vdd.n503 361.584
R2288 vdd.n567 vdd.n534 361.584
R2289 vdd.n718 vdd.n717 361.584
R2290 vdd.n758 vdd.n448 361.584
R2291 vdd.n774 vdd.n773 361.584
R2292 vdd.n645 vdd.n578 349.733
R2293 vdd.n781 vdd.n47 349.733
R2294 vdd.n817 vdd.n11 349.733
R2295 vdd.n638 vdd.n637 341.769
R2296 vdd.n68 vdd.n46 341.769
R2297 vdd.n795 vdd.n29 341.769
R2298 vdd.n789 vdd.n788 304.478
R2299 vdd.n32 vdd.n31 294.932
R2300 vdd.n583 vdd.n581 285.291
R2301 vdd.n75 vdd.n38 285.291
R2302 vdd.n626 vdd.n625 269.361
R2303 vdd.n60 vdd.n56 269.361
R2304 vdd.n790 vdd.n28 269.361
R2305 vdd.n19 vdd.n14 245.827
R2306 vdd.n10 vdd.n8 201.326
R2307 vdd.n622 vdd.n619 190.871
R2308 vdd.n619 vdd.n617 190.871
R2309 vdd.n432 vdd 190.871
R2310 vdd.n409 vdd 190.871
R2311 vdd.n432 vdd.n431 190.871
R2312 vdd.n405 vdd 190.871
R2313 vdd.n436 vdd 190.871
R2314 vdd.n405 vdd.n399 190.871
R2315 vdd.n415 vdd.n410 190.871
R2316 vdd.n415 vdd 190.871
R2317 vdd.n426 vdd 190.871
R2318 vdd.n422 vdd 190.871
R2319 vdd vdd.n421 190.871
R2320 vdd.n421 vdd.n420 190.871
R2321 vdd.n152 vdd.n143 190.871
R2322 vdd.n152 vdd 190.871
R2323 vdd vdd.n151 190.871
R2324 vdd.n158 vdd.n138 190.871
R2325 vdd.n158 vdd 190.871
R2326 vdd vdd.n157 190.871
R2327 vdd.n125 vdd.n124 190.871
R2328 vdd.n124 vdd 190.871
R2329 vdd.n164 vdd.n85 190.871
R2330 vdd vdd.n85 190.871
R2331 vdd.n117 vdd.n100 190.871
R2332 vdd vdd.n117 190.871
R2333 vdd.n118 vdd 190.871
R2334 vdd.n112 vdd 190.871
R2335 vdd vdd.n111 190.871
R2336 vdd.n111 vdd.n108 190.871
R2337 vdd.n548 vdd.n502 190.871
R2338 vdd.n548 vdd.n547 190.871
R2339 vdd.n715 vdd.n695 190.871
R2340 vdd.n695 vdd.n694 190.871
R2341 vdd.n702 vdd.n480 190.871
R2342 vdd.n703 vdd.n702 190.871
R2343 vdd.n529 vdd.n492 190.871
R2344 vdd.n686 vdd.n492 190.871
R2345 vdd.n783 vdd.n43 190.871
R2346 vdd.n784 vdd.n783 190.871
R2347 vdd.n813 vdd.n812 190.871
R2348 vdd.n812 vdd.n25 190.871
R2349 vdd.n202 vdd 190.871
R2350 vdd.n211 vdd 190.871
R2351 vdd.n202 vdd.n187 190.871
R2352 vdd.n218 vdd 190.871
R2353 vdd.n183 vdd 190.871
R2354 vdd.n218 vdd.n217 190.871
R2355 vdd vdd.n330 190.871
R2356 vdd.n330 vdd.n329 190.871
R2357 vdd vdd.n174 190.871
R2358 vdd.n346 vdd.n174 190.871
R2359 vdd.n304 vdd 190.871
R2360 vdd.n304 vdd.n303 190.871
R2361 vdd.n318 vdd 190.871
R2362 vdd.n318 vdd.n317 190.871
R2363 vdd.n278 vdd 190.871
R2364 vdd.n309 vdd 190.871
R2365 vdd.n278 vdd.n250 190.871
R2366 vdd.n270 vdd 190.871
R2367 vdd.n265 vdd 190.871
R2368 vdd.n270 vdd.n269 190.871
R2369 vdd.n206 vdd.n193 190.871
R2370 vdd vdd.n206 190.871
R2371 vdd.n207 vdd 190.871
R2372 vdd.n197 vdd.n196 190.871
R2373 vdd vdd.n197 190.871
R2374 vdd.n198 vdd 190.871
R2375 vdd.n243 vdd.n232 190.871
R2376 vdd vdd.n243 190.871
R2377 vdd.n239 vdd.n237 190.871
R2378 vdd vdd.n239 190.871
R2379 vdd.n282 vdd.n256 190.871
R2380 vdd vdd.n282 190.871
R2381 vdd.n283 vdd 190.871
R2382 vdd.n275 vdd 190.871
R2383 vdd vdd.n274 190.871
R2384 vdd.n274 vdd.n262 190.871
R2385 vdd.n388 vdd 190.871
R2386 vdd.n365 vdd 190.871
R2387 vdd.n388 vdd.n387 190.871
R2388 vdd.n361 vdd 190.871
R2389 vdd.n392 vdd 190.871
R2390 vdd.n361 vdd.n355 190.871
R2391 vdd.n371 vdd.n366 190.871
R2392 vdd.n371 vdd 190.871
R2393 vdd.n382 vdd 190.871
R2394 vdd.n378 vdd 190.871
R2395 vdd vdd.n377 190.871
R2396 vdd.n377 vdd.n376 190.871
R2397 vdd.n430 vdd.n409 190.494
R2398 vdd.n437 vdd.n436 190.494
R2399 vdd.n427 vdd.n426 190.494
R2400 vdd.n422 vdd.n397 190.494
R2401 vdd.n151 vdd.n148 190.494
R2402 vdd.n157 vdd.n139 190.494
R2403 vdd.n118 vdd.n99 190.494
R2404 vdd.n112 vdd.n107 190.494
R2405 vdd.n212 vdd.n211 190.494
R2406 vdd.n216 vdd.n183 190.494
R2407 vdd.n310 vdd.n309 190.494
R2408 vdd.n268 vdd.n265 190.494
R2409 vdd.n207 vdd.n185 190.494
R2410 vdd.n198 vdd.n184 190.494
R2411 vdd.n283 vdd.n249 190.494
R2412 vdd.n275 vdd.n261 190.494
R2413 vdd.n386 vdd.n365 190.494
R2414 vdd.n393 vdd.n392 190.494
R2415 vdd.n383 vdd.n382 190.494
R2416 vdd.n378 vdd.n353 190.494
R2417 vdd.n20 vdd.n10 185
R2418 vdd.n114 vdd.n101 179.118
R2419 vdd.n115 vdd.n96 179.118
R2420 vdd.n120 vdd.n96 179.118
R2421 vdd.n122 vdd.n121 179.118
R2422 vdd.n121 vdd.n93 179.118
R2423 vdd.n131 vdd.n93 179.118
R2424 vdd.n131 vdd.n88 179.118
R2425 vdd.n162 vdd.n88 179.118
R2426 vdd.n162 vdd.n161 179.118
R2427 vdd.n160 vdd.n135 179.118
R2428 vdd.n155 vdd.n135 179.118
R2429 vdd.n154 vdd.n140 179.118
R2430 vdd.n756 vdd.n451 174.868
R2431 vdd.n512 vdd.n496 174.868
R2432 vdd.n110 vdd.n109 173.642
R2433 vdd.n150 vdd.n149 173.642
R2434 vdd.n748 vdd.n464 170.885
R2435 vdd.n675 vdd.n508 170.885
R2436 vdd.n727 vdd.n690 152.239
R2437 vdd.n721 vdd.n486 142.645
R2438 vdd.n666 vdd.n499 142.645
R2439 vdd.n20 vdd.n16 137.326
R2440 vdd.n627 vdd.n626 136.964
R2441 vdd.n60 vdd.n55 136.964
R2442 vdd.n742 vdd.n471 134.68
R2443 vdd.n543 vdd.n488 134.68
R2444 vdd.n165 vdd.n84 131.388
R2445 vdd.n133 vdd.n84 131.388
R2446 vdd.n127 vdd.n126 131.388
R2447 vdd.n127 vdd.n91 131.388
R2448 vdd.n342 vdd.n173 131.388
R2449 vdd.n347 vdd.n173 131.388
R2450 vdd.n327 vdd.n225 131.388
R2451 vdd.n328 vdd.n327 131.388
R2452 vdd.n296 vdd.n247 131.388
R2453 vdd.n316 vdd.n247 131.388
R2454 vdd.n301 vdd.n288 131.388
R2455 vdd.n302 vdd.n301 131.388
R2456 vdd.n236 vdd.n235 131.388
R2457 vdd.n240 vdd.n235 131.388
R2458 vdd.n337 vdd.n336 131.388
R2459 vdd.n336 vdd.n241 131.388
R2460 vdd.n21 vdd.n20 123.334
R2461 vdd.n599 vdd.n583 123.096
R2462 vdd.n788 vdd.n38 123.096
R2463 vdd.n790 vdd.n789 122.733
R2464 vdd.n161 vdd.n160 120.168
R2465 vdd.n115 vdd.n114 117.9
R2466 vdd.n155 vdd.n154 117.9
R2467 vdd.n793 vdd.n17 98.5799
R2468 vdd.n412 vdd 92.5005
R2469 vdd.n417 vdd.n412 92.5005
R2470 vdd.n411 vdd.n410 92.5005
R2471 vdd.n413 vdd.n411 92.5005
R2472 vdd.n401 vdd.n399 92.5005
R2473 vdd.n404 vdd.n401 92.5005
R2474 vdd.n400 vdd 92.5005
R2475 vdd.n402 vdd.n400 92.5005
R2476 vdd.n431 vdd.n408 92.5005
R2477 vdd.n408 vdd.n404 92.5005
R2478 vdd vdd.n407 92.5005
R2479 vdd.n407 vdd.n402 92.5005
R2480 vdd vdd.n419 92.5005
R2481 vdd.n419 vdd.n417 92.5005
R2482 vdd.n420 vdd.n418 92.5005
R2483 vdd.n418 vdd.n413 92.5005
R2484 vdd vdd.n98 92.5005
R2485 vdd.n98 vdd.n96 92.5005
R2486 vdd.n100 vdd.n97 92.5005
R2487 vdd.n97 vdd.n96 92.5005
R2488 vdd.n134 vdd 92.5005
R2489 vdd.n162 vdd.n134 92.5005
R2490 vdd vdd.n132 92.5005
R2491 vdd.n132 vdd.n131 92.5005
R2492 vdd.n95 vdd 92.5005
R2493 vdd.n121 vdd.n95 92.5005
R2494 vdd.n125 vdd.n94 92.5005
R2495 vdd.n121 vdd.n94 92.5005
R2496 vdd.n130 vdd.n83 92.5005
R2497 vdd.n131 vdd.n130 92.5005
R2498 vdd.n164 vdd.n163 92.5005
R2499 vdd.n163 vdd.n162 92.5005
R2500 vdd vdd.n137 92.5005
R2501 vdd.n137 vdd.n135 92.5005
R2502 vdd.n138 vdd.n136 92.5005
R2503 vdd.n136 vdd.n135 92.5005
R2504 vdd vdd.n142 92.5005
R2505 vdd.n143 vdd.n141 92.5005
R2506 vdd.n141 vdd.n140 92.5005
R2507 vdd vdd.n103 92.5005
R2508 vdd.n103 vdd.n101 92.5005
R2509 vdd.n108 vdd.n102 92.5005
R2510 vdd vdd.n255 92.5005
R2511 vdd.n255 vdd.n253 92.5005
R2512 vdd.n256 vdd.n254 92.5005
R2513 vdd.n254 vdd.n253 92.5005
R2514 vdd vdd.n178 92.5005
R2515 vdd.n344 vdd.n178 92.5005
R2516 vdd vdd.n229 92.5005
R2517 vdd.n340 vdd.n229 92.5005
R2518 vdd.n333 vdd 92.5005
R2519 vdd.n333 vdd.n332 92.5005
R2520 vdd.n323 vdd.n232 92.5005
R2521 vdd.n332 vdd.n323 92.5005
R2522 vdd.n339 vdd.n338 92.5005
R2523 vdd.n340 vdd.n339 92.5005
R2524 vdd.n237 vdd.n222 92.5005
R2525 vdd.n344 vdd.n222 92.5005
R2526 vdd vdd.n195 92.5005
R2527 vdd.n195 vdd.n180 92.5005
R2528 vdd.n196 vdd.n194 92.5005
R2529 vdd.n194 vdd.n180 92.5005
R2530 vdd vdd.n192 92.5005
R2531 vdd.n192 vdd.n190 92.5005
R2532 vdd.n193 vdd.n191 92.5005
R2533 vdd.n191 vdd.n190 92.5005
R2534 vdd.n269 vdd.n264 92.5005
R2535 vdd.n264 vdd.n257 92.5005
R2536 vdd vdd.n263 92.5005
R2537 vdd.n263 vdd.n257 92.5005
R2538 vdd.n252 vdd.n250 92.5005
R2539 vdd.n253 vdd.n252 92.5005
R2540 vdd.n251 vdd 92.5005
R2541 vdd.n253 vdd.n251 92.5005
R2542 vdd.n317 vdd.n246 92.5005
R2543 vdd.n246 vdd.n244 92.5005
R2544 vdd.n291 vdd.n248 92.5005
R2545 vdd.n298 vdd.n291 92.5005
R2546 vdd.n303 vdd.n287 92.5005
R2547 vdd.n287 vdd.n285 92.5005
R2548 vdd vdd.n286 92.5005
R2549 vdd.n286 vdd.n285 92.5005
R2550 vdd.n297 vdd 92.5005
R2551 vdd.n298 vdd.n297 92.5005
R2552 vdd vdd.n245 92.5005
R2553 vdd.n245 vdd.n244 92.5005
R2554 vdd.n346 vdd.n345 92.5005
R2555 vdd.n345 vdd.n344 92.5005
R2556 vdd.n228 vdd.n172 92.5005
R2557 vdd.n340 vdd.n228 92.5005
R2558 vdd.n329 vdd.n322 92.5005
R2559 vdd.n332 vdd.n322 92.5005
R2560 vdd.n331 vdd 92.5005
R2561 vdd.n332 vdd.n331 92.5005
R2562 vdd vdd.n341 92.5005
R2563 vdd.n341 vdd.n340 92.5005
R2564 vdd.n343 vdd 92.5005
R2565 vdd.n344 vdd.n343 92.5005
R2566 vdd.n217 vdd.n182 92.5005
R2567 vdd.n182 vdd.n180 92.5005
R2568 vdd vdd.n181 92.5005
R2569 vdd.n181 vdd.n180 92.5005
R2570 vdd.n189 vdd.n187 92.5005
R2571 vdd.n190 vdd.n189 92.5005
R2572 vdd.n188 vdd 92.5005
R2573 vdd.n190 vdd.n188 92.5005
R2574 vdd vdd.n260 92.5005
R2575 vdd.n260 vdd.n257 92.5005
R2576 vdd.n262 vdd.n259 92.5005
R2577 vdd.n259 vdd.n257 92.5005
R2578 vdd.n368 vdd 92.5005
R2579 vdd.n373 vdd.n368 92.5005
R2580 vdd.n367 vdd.n366 92.5005
R2581 vdd.n369 vdd.n367 92.5005
R2582 vdd.n357 vdd.n355 92.5005
R2583 vdd.n360 vdd.n357 92.5005
R2584 vdd.n356 vdd 92.5005
R2585 vdd.n358 vdd.n356 92.5005
R2586 vdd.n387 vdd.n364 92.5005
R2587 vdd.n364 vdd.n360 92.5005
R2588 vdd vdd.n363 92.5005
R2589 vdd.n363 vdd.n358 92.5005
R2590 vdd vdd.n375 92.5005
R2591 vdd.n375 vdd.n373 92.5005
R2592 vdd.n376 vdd.n374 92.5005
R2593 vdd.n374 vdd.n369 92.5005
R2594 vdd.n434 vdd.n402 91.6935
R2595 vdd.n434 vdd.n404 91.6935
R2596 vdd.n424 vdd.n413 91.6935
R2597 vdd.n424 vdd.n417 91.6935
R2598 vdd.n390 vdd.n358 91.6935
R2599 vdd.n390 vdd.n360 91.6935
R2600 vdd.n380 vdd.n369 91.6935
R2601 vdd.n380 vdd.n373 91.6935
R2602 vdd.n272 vdd.n257 89.559
R2603 vdd.n277 vdd.n257 89.559
R2604 vdd.n280 vdd.n253 89.559
R2605 vdd.n307 vdd.n253 89.559
R2606 vdd.n306 vdd.n285 89.559
R2607 vdd.n299 vdd.n285 89.559
R2608 vdd.n299 vdd.n298 89.559
R2609 vdd.n298 vdd.n292 89.559
R2610 vdd.n292 vdd.n244 89.559
R2611 vdd.n320 vdd.n244 89.559
R2612 vdd.n332 vdd.n321 89.559
R2613 vdd.n332 vdd.n227 89.559
R2614 vdd.n340 vdd.n227 89.559
R2615 vdd.n340 vdd.n177 89.559
R2616 vdd.n344 vdd.n177 89.559
R2617 vdd.n344 vdd.n221 89.559
R2618 vdd.n220 vdd.n180 89.559
R2619 vdd.n201 vdd.n180 89.559
R2620 vdd.n204 vdd.n190 89.559
R2621 vdd.n209 vdd.n190 89.559
R2622 vdd.n609 vdd.n608 85.0829
R2623 vdd.n609 vdd.n574 85.0829
R2624 vdd.n564 vdd.n539 85.0829
R2625 vdd.n565 vdd.n564 85.0829
R2626 vdd.n753 vdd.n752 85.0829
R2627 vdd.n752 vdd.n459 85.0829
R2628 vdd.n735 vdd.n447 85.0829
R2629 vdd.n736 vdd.n735 85.0829
R2630 vdd.n671 vdd.n517 85.0829
R2631 vdd.n672 vdd.n671 85.0829
R2632 vdd.n779 vdd.n50 85.0829
R2633 vdd.n779 vdd.n778 85.0829
R2634 vdd.n800 vdd.n7 85.0829
R2635 vdd.n800 vdd.n799 85.0829
R2636 vdd.n149 vdd.n142 79.4196
R2637 vdd.n109 vdd.n102 79.4196
R2638 vdd.n617 vdd.n601 66.7857
R2639 vdd.n547 vdd.n546 66.7857
R2640 vdd.n694 vdd.n457 66.7857
R2641 vdd.n731 vdd.n480 66.7857
R2642 vdd.n530 vdd.n529 66.7857
R2643 vdd.n79 vdd.n43 66.7857
R2644 vdd.n814 vdd.n813 66.7857
R2645 vdd.n814 vdd.n17 66.6358
R2646 vdd.n629 vdd.n615 66.1931
R2647 vdd.n544 vdd.n542 66.1931
R2648 vdd.n693 vdd.n466 66.1931
R2649 vdd.n479 vdd.n478 66.1931
R2650 vdd.n528 vdd.n527 66.1931
R2651 vdd.n72 vdd.n71 66.1931
R2652 vdd.n806 vdd.n18 66.1931
R2653 vdd.n637 vdd.n606 62.6339
R2654 vdd.n69 vdd.n68 62.6339
R2655 vdd.n808 vdd.n29 62.6339
R2656 vdd.n727 vdd.n486 61.5478
R2657 vdd.n666 vdd.n535 61.5478
R2658 vdd.n707 vdd.n471 61.3667
R2659 vdd.n690 vdd.n488 61.3667
R2660 vdd.n645 vdd.n644 60.4616
R2661 vdd.n74 vdd.n47 60.4616
R2662 vdd.n817 vdd.n816 60.4616
R2663 vdd.n307 vdd.n306 60.084
R2664 vdd.n321 vdd.n320 60.084
R2665 vdd.n221 vdd.n220 60.084
R2666 vdd.n126 vdd.n125 59.4829
R2667 vdd.n126 vdd.n83 59.4829
R2668 vdd.n165 vdd.n164 59.4829
R2669 vdd vdd.n91 59.4829
R2670 vdd vdd.n91 59.4829
R2671 vdd.n133 vdd 59.4829
R2672 vdd vdd.n133 59.4829
R2673 vdd vdd.n225 59.4829
R2674 vdd vdd.n225 59.4829
R2675 vdd.n342 vdd 59.4829
R2676 vdd vdd.n342 59.4829
R2677 vdd.n329 vdd.n328 59.4829
R2678 vdd.n328 vdd.n172 59.4829
R2679 vdd.n347 vdd.n346 59.4829
R2680 vdd.n288 vdd 59.4829
R2681 vdd vdd.n288 59.4829
R2682 vdd vdd.n296 59.4829
R2683 vdd.n296 vdd 59.4829
R2684 vdd.n303 vdd.n302 59.4829
R2685 vdd.n302 vdd.n248 59.4829
R2686 vdd.n317 vdd.n316 59.4829
R2687 vdd.n337 vdd.n232 59.4829
R2688 vdd.n338 vdd.n337 59.4829
R2689 vdd.n237 vdd.n236 59.4829
R2690 vdd vdd.n241 59.4829
R2691 vdd.n241 vdd 59.4829
R2692 vdd vdd.n240 59.4829
R2693 vdd.n240 vdd 59.4829
R2694 vdd.n166 vdd.n165 59.1064
R2695 vdd.n348 vdd.n347 59.1064
R2696 vdd.n316 vdd.n315 59.1064
R2697 vdd.n236 vdd.n170 59.1064
R2698 vdd.n280 vdd.n277 58.9504
R2699 vdd.n204 vdd.n201 58.9504
R2700 vdd.n799 vdd.n798 53.6992
R2701 vdd.n608 vdd.n607 52.3937
R2702 vdd.n545 vdd.n539 52.3937
R2703 vdd.n754 vdd.n753 52.3937
R2704 vdd.n736 vdd.n732 52.3937
R2705 vdd.n672 vdd.n516 52.3937
R2706 vdd.n778 vdd.n777 52.3937
R2707 vdd.n630 vdd.n605 51.2005
R2708 vdd.n560 vdd.n507 51.2005
R2709 vdd.n746 vdd.n458 51.2005
R2710 vdd.n738 vdd.n737 51.2005
R2711 vdd.n673 vdd.n515 51.2005
R2712 vdd.n58 vdd.n51 51.2005
R2713 vdd.n804 vdd.n32 48.9418
R2714 vdd.n793 vdd.n14 46.2505
R2715 vdd.n815 vdd.n814 40.0406
R2716 vdd.n20 vdd.n19 39.4632
R2717 vdd vdd.n589 37.0005
R2718 vdd.n597 vdd.n596 37.0005
R2719 vdd.n598 vdd.n597 37.0005
R2720 vdd.n641 vdd.n640 37.0005
R2721 vdd.n640 vdd.n581 37.0005
R2722 vdd.n577 vdd.n575 37.0005
R2723 vdd.n583 vdd.n577 37.0005
R2724 vdd.n634 vdd.n613 37.0005
R2725 vdd.n626 vdd.n613 37.0005
R2726 vdd.n632 vdd.n604 37.0005
R2727 vdd.n625 vdd.n604 37.0005
R2728 vdd.n610 vdd.n609 37.0005
R2729 vdd.n610 vdd.n578 37.0005
R2730 vdd.n720 vdd.n481 37.0005
R2731 vdd.n721 vdd.n720 37.0005
R2732 vdd.n741 vdd.n740 37.0005
R2733 vdd.n742 vdd.n741 37.0005
R2734 vdd.n735 vdd.n734 37.0005
R2735 vdd.n734 vdd.n451 37.0005
R2736 vdd.n450 vdd.n448 37.0005
R2737 vdd.n486 vdd.n450 37.0005
R2738 vdd.n476 vdd.n475 37.0005
R2739 vdd.n475 vdd.n471 37.0005
R2740 vdd.n667 vdd.n534 37.0005
R2741 vdd.n667 vdd.n666 37.0005
R2742 vdd.n522 vdd.n521 37.0005
R2743 vdd.n522 vdd.n488 37.0005
R2744 vdd.n752 vdd.n751 37.0005
R2745 vdd.n751 vdd.n451 37.0005
R2746 vdd.n718 vdd.n456 37.0005
R2747 vdd.n486 vdd.n456 37.0005
R2748 vdd.n467 vdd.n460 37.0005
R2749 vdd.n471 vdd.n460 37.0005
R2750 vdd.n564 vdd.n563 37.0005
R2751 vdd.n563 vdd.n512 37.0005
R2752 vdd.n665 vdd.n503 37.0005
R2753 vdd.n666 vdd.n665 37.0005
R2754 vdd.n556 vdd.n541 37.0005
R2755 vdd.n541 vdd.n488 37.0005
R2756 vdd.n723 vdd.n722 37.0005
R2757 vdd.n722 vdd.n721 37.0005
R2758 vdd.n744 vdd.n743 37.0005
R2759 vdd.n743 vdd.n742 37.0005
R2760 vdd.n678 vdd.n677 37.0005
R2761 vdd.n677 vdd.n499 37.0005
R2762 vdd.n558 vdd.n506 37.0005
R2763 vdd.n543 vdd.n506 37.0005
R2764 vdd.n532 vdd.n514 37.0005
R2765 vdd.n514 vdd.n499 37.0005
R2766 vdd.n525 vdd.n513 37.0005
R2767 vdd.n543 vdd.n513 37.0005
R2768 vdd.n671 vdd.n670 37.0005
R2769 vdd.n670 vdd.n512 37.0005
R2770 vdd.n77 vdd.n76 37.0005
R2771 vdd.n76 vdd.n75 37.0005
R2772 vdd.n63 vdd.n53 37.0005
R2773 vdd.n56 vdd.n53 37.0005
R2774 vdd.n780 vdd.n779 37.0005
R2775 vdd.n781 vdd.n780 37.0005
R2776 vdd.n775 vdd.n774 37.0005
R2777 vdd.n775 vdd.n38 37.0005
R2778 vdd.n65 vdd.n61 37.0005
R2779 vdd.n61 vdd.n60 37.0005
R2780 vdd.n791 vdd.n37 37.0005
R2781 vdd.n791 vdd.n790 37.0005
R2782 vdd.n792 vdd.n30 37.0005
R2783 vdd.n792 vdd.n28 37.0005
R2784 vdd.n801 vdd.n800 37.0005
R2785 vdd.n801 vdd.n11 37.0005
R2786 vdd.n23 vdd.n22 32.7398
R2787 vdd.n748 vdd.n462 31.3172
R2788 vdd.n552 vdd.n508 31.3172
R2789 vdd.n756 vdd.n454 30.2311
R2790 vdd.n683 vdd.n496 30.2311
R2791 vdd.n633 vdd.n614 26.6787
R2792 vdd.n557 vdd.n555 26.6787
R2793 vdd.n696 vdd.n468 26.6787
R2794 vdd.n705 vdd.n477 26.6787
R2795 vdd.n688 vdd.n491 26.6787
R2796 vdd.n64 vdd.n62 26.6787
R2797 vdd.n36 vdd.n35 26.6787
R2798 vdd.n620 vdd.n602 26.63
R2799 vdd.n680 vdd.n679 26.63
R2800 vdd.n725 vdd.n724 26.63
R2801 vdd.n485 vdd.n484 26.63
R2802 vdd.n533 vdd.n493 26.63
R2803 vdd.n786 vdd.n41 26.63
R2804 vdd.n413 vdd.n404 26.5564
R2805 vdd.n369 vdd.n360 26.5564
R2806 vdd.n426 vdd.n425 23.1255
R2807 vdd.n425 vdd.n424 23.1255
R2808 vdd.n416 vdd.n415 23.1255
R2809 vdd.n424 vdd.n416 23.1255
R2810 vdd.n436 vdd.n435 23.1255
R2811 vdd.n435 vdd.n434 23.1255
R2812 vdd.n406 vdd.n405 23.1255
R2813 vdd.n434 vdd.n406 23.1255
R2814 vdd.n409 vdd.n403 23.1255
R2815 vdd.n434 vdd.n403 23.1255
R2816 vdd.n433 vdd.n432 23.1255
R2817 vdd.n434 vdd.n433 23.1255
R2818 vdd.n423 vdd.n422 23.1255
R2819 vdd.n424 vdd.n423 23.1255
R2820 vdd.n421 vdd.n414 23.1255
R2821 vdd.n424 vdd.n414 23.1255
R2822 vdd.n119 vdd.n118 23.1255
R2823 vdd.n120 vdd.n119 23.1255
R2824 vdd.n117 vdd.n116 23.1255
R2825 vdd.n116 vdd.n115 23.1255
R2826 vdd.n128 vdd.n127 23.1255
R2827 vdd.n128 vdd.n93 23.1255
R2828 vdd.n89 vdd.n84 23.1255
R2829 vdd.n89 vdd.n88 23.1255
R2830 vdd.n87 vdd.n85 23.1255
R2831 vdd.n161 vdd.n87 23.1255
R2832 vdd.n124 vdd.n123 23.1255
R2833 vdd.n123 vdd.n122 23.1255
R2834 vdd.n157 vdd.n156 23.1255
R2835 vdd.n156 vdd.n155 23.1255
R2836 vdd.n159 vdd.n158 23.1255
R2837 vdd.n160 vdd.n159 23.1255
R2838 vdd.n151 vdd.n150 23.1255
R2839 vdd.n153 vdd.n152 23.1255
R2840 vdd.n154 vdd.n153 23.1255
R2841 vdd.n113 vdd.n112 23.1255
R2842 vdd.n114 vdd.n113 23.1255
R2843 vdd.n111 vdd.n110 23.1255
R2844 vdd.n284 vdd.n283 23.1255
R2845 vdd.n307 vdd.n284 23.1255
R2846 vdd.n282 vdd.n281 23.1255
R2847 vdd.n281 vdd.n280 23.1255
R2848 vdd.n336 vdd.n335 23.1255
R2849 vdd.n335 vdd.n227 23.1255
R2850 vdd.n235 vdd.n234 23.1255
R2851 vdd.n234 vdd.n177 23.1255
R2852 vdd.n239 vdd.n238 23.1255
R2853 vdd.n238 vdd.n221 23.1255
R2854 vdd.n243 vdd.n242 23.1255
R2855 vdd.n321 vdd.n242 23.1255
R2856 vdd.n199 vdd.n198 23.1255
R2857 vdd.n201 vdd.n199 23.1255
R2858 vdd.n197 vdd.n179 23.1255
R2859 vdd.n220 vdd.n179 23.1255
R2860 vdd.n208 vdd.n207 23.1255
R2861 vdd.n209 vdd.n208 23.1255
R2862 vdd.n206 vdd.n205 23.1255
R2863 vdd.n205 vdd.n204 23.1255
R2864 vdd.n265 vdd.n258 23.1255
R2865 vdd.n277 vdd.n258 23.1255
R2866 vdd.n271 vdd.n270 23.1255
R2867 vdd.n272 vdd.n271 23.1255
R2868 vdd.n309 vdd.n308 23.1255
R2869 vdd.n308 vdd.n307 23.1255
R2870 vdd.n279 vdd.n278 23.1255
R2871 vdd.n280 vdd.n279 23.1255
R2872 vdd.n301 vdd.n300 23.1255
R2873 vdd.n300 vdd.n299 23.1255
R2874 vdd.n294 vdd.n247 23.1255
R2875 vdd.n294 vdd.n292 23.1255
R2876 vdd.n319 vdd.n318 23.1255
R2877 vdd.n320 vdd.n319 23.1255
R2878 vdd.n305 vdd.n304 23.1255
R2879 vdd.n306 vdd.n305 23.1255
R2880 vdd.n327 vdd.n326 23.1255
R2881 vdd.n326 vdd.n227 23.1255
R2882 vdd.n223 vdd.n173 23.1255
R2883 vdd.n223 vdd.n177 23.1255
R2884 vdd.n176 vdd.n174 23.1255
R2885 vdd.n221 vdd.n176 23.1255
R2886 vdd.n330 vdd.n324 23.1255
R2887 vdd.n324 vdd.n321 23.1255
R2888 vdd.n200 vdd.n183 23.1255
R2889 vdd.n201 vdd.n200 23.1255
R2890 vdd.n219 vdd.n218 23.1255
R2891 vdd.n220 vdd.n219 23.1255
R2892 vdd.n211 vdd.n210 23.1255
R2893 vdd.n210 vdd.n209 23.1255
R2894 vdd.n203 vdd.n202 23.1255
R2895 vdd.n204 vdd.n203 23.1255
R2896 vdd.n276 vdd.n275 23.1255
R2897 vdd.n277 vdd.n276 23.1255
R2898 vdd.n274 vdd.n273 23.1255
R2899 vdd.n273 vdd.n272 23.1255
R2900 vdd.n382 vdd.n381 23.1255
R2901 vdd.n381 vdd.n380 23.1255
R2902 vdd.n372 vdd.n371 23.1255
R2903 vdd.n380 vdd.n372 23.1255
R2904 vdd.n392 vdd.n391 23.1255
R2905 vdd.n391 vdd.n390 23.1255
R2906 vdd.n362 vdd.n361 23.1255
R2907 vdd.n390 vdd.n362 23.1255
R2908 vdd.n365 vdd.n359 23.1255
R2909 vdd.n390 vdd.n359 23.1255
R2910 vdd.n389 vdd.n388 23.1255
R2911 vdd.n390 vdd.n389 23.1255
R2912 vdd.n379 vdd.n378 23.1255
R2913 vdd.n380 vdd.n379 23.1255
R2914 vdd.n377 vdd.n370 23.1255
R2915 vdd.n380 vdd.n370 23.1255
R2916 vdd.n798 vdd.n17 19.2575
R2917 vdd.n631 vdd.n630 19.0689
R2918 vdd.n560 vdd.n559 19.0689
R2919 vdd.n746 vdd.n745 19.0689
R2920 vdd.n739 vdd.n738 19.0689
R2921 vdd.n526 vdd.n515 19.0689
R2922 vdd.n58 vdd.n54 19.0689
R2923 vdd.n805 vdd.n804 19.0689
R2924 vdd.n625 vdd.n606 17.7406
R2925 vdd.n69 vdd.n56 17.7406
R2926 vdd.n808 vdd.n28 17.7406
R2927 vdd.n641 vdd.n602 17.4344
R2928 vdd.n679 vdd.n678 17.4344
R2929 vdd.n724 vdd.n723 17.4344
R2930 vdd.n484 vdd.n481 17.4344
R2931 vdd.n533 vdd.n532 17.4344
R2932 vdd.n77 vdd.n41 17.4344
R2933 vdd.n607 vdd.n601 16.8923
R2934 vdd.n530 vdd.n516 16.8923
R2935 vdd.n546 vdd.n545 16.8923
R2936 vdd.n754 vdd.n457 16.8923
R2937 vdd.n732 vdd.n731 16.8923
R2938 vdd.n777 vdd.n79 16.8923
R2939 vdd.n633 vdd.n632 16.6793
R2940 vdd.n558 vdd.n557 16.6793
R2941 vdd.n744 vdd.n468 16.6793
R2942 vdd.n740 vdd.n477 16.6793
R2943 vdd.n525 vdd.n491 16.6793
R2944 vdd.n64 vdd.n63 16.6793
R2945 vdd.n36 vdd.n30 16.6793
R2946 vdd.n627 vdd.n614 14.2313
R2947 vdd.n619 vdd.n618 14.2313
R2948 vdd.n618 vdd.n578 14.2313
R2949 vdd.n620 vdd.n600 14.2313
R2950 vdd.n600 vdd.n599 14.2313
R2951 vdd.n702 vdd.n701 14.2313
R2952 vdd.n701 vdd.n451 14.2313
R2953 vdd.n728 vdd.n485 14.2313
R2954 vdd.n728 vdd.n727 14.2313
R2955 vdd.n706 vdd.n705 14.2313
R2956 vdd.n707 vdd.n706 14.2313
R2957 vdd.n711 vdd.n695 14.2313
R2958 vdd.n711 vdd.n451 14.2313
R2959 vdd.n726 vdd.n725 14.2313
R2960 vdd.n727 vdd.n726 14.2313
R2961 vdd.n708 vdd.n696 14.2313
R2962 vdd.n708 vdd.n707 14.2313
R2963 vdd.n549 vdd.n548 14.2313
R2964 vdd.n549 vdd.n512 14.2313
R2965 vdd.n680 vdd.n501 14.2313
R2966 vdd.n535 vdd.n501 14.2313
R2967 vdd.n555 vdd.n487 14.2313
R2968 vdd.n690 vdd.n487 14.2313
R2969 vdd.n495 vdd.n493 14.2313
R2970 vdd.n535 vdd.n495 14.2313
R2971 vdd.n511 vdd.n492 14.2313
R2972 vdd.n512 vdd.n511 14.2313
R2973 vdd.n689 vdd.n688 14.2313
R2974 vdd.n690 vdd.n689 14.2313
R2975 vdd.n783 vdd.n782 14.2313
R2976 vdd.n782 vdd.n781 14.2313
R2977 vdd.n787 vdd.n786 14.2313
R2978 vdd.n788 vdd.n787 14.2313
R2979 vdd.n62 vdd.n55 14.2313
R2980 vdd.n23 vdd.n16 14.2313
R2981 vdd.n812 vdd.n811 14.2313
R2982 vdd.n811 vdd.n11 14.2313
R2983 vdd.n35 vdd.n26 14.2313
R2984 vdd.n789 vdd.n26 14.2313
R2985 vdd.n22 vdd.n17 12.6319
R2986 vdd.n149 vdd.n140 8.97701
R2987 vdd.n109 vdd.n101 8.97701
R2988 vdd.n742 vdd.n462 8.87055
R2989 vdd.n552 vdd.n543 8.87055
R2990 vdd.n22 vdd.n21 8.1562
R2991 vdd.n638 vdd.n578 7.96544
R2992 vdd.n781 vdd.n46 7.96544
R2993 vdd.n795 vdd.n11 7.96544
R2994 vdd.n630 vdd.n612 7.11588
R2995 vdd.n637 vdd.n612 7.11588
R2996 vdd.n607 vdd.n579 7.11588
R2997 vdd.n645 vdd.n579 7.11588
R2998 vdd.n647 vdd.n646 7.11588
R2999 vdd.n646 vdd.n645 7.11588
R3000 vdd.n636 vdd.n635 7.11588
R3001 vdd.n637 vdd.n636 7.11588
R3002 vdd.n732 vdd.n453 7.11588
R3003 vdd.n756 vdd.n453 7.11588
R3004 vdd.n738 vdd.n463 7.11588
R3005 vdd.n748 vdd.n463 7.11588
R3006 vdd.n474 vdd.n465 7.11588
R3007 vdd.n748 vdd.n465 7.11588
R3008 vdd.n758 vdd.n757 7.11588
R3009 vdd.n757 vdd.n756 7.11588
R3010 vdd.n717 vdd.n452 7.11588
R3011 vdd.n756 vdd.n452 7.11588
R3012 vdd.n749 vdd.n461 7.11588
R3013 vdd.n749 vdd.n748 7.11588
R3014 vdd.n747 vdd.n746 7.11588
R3015 vdd.n748 vdd.n747 7.11588
R3016 vdd.n755 vdd.n754 7.11588
R3017 vdd.n756 vdd.n755 7.11588
R3018 vdd.n664 vdd.n663 7.11588
R3019 vdd.n664 vdd.n496 7.11588
R3020 vdd.n540 vdd.n538 7.11588
R3021 vdd.n540 vdd.n508 7.11588
R3022 vdd.n561 vdd.n560 7.11588
R3023 vdd.n561 vdd.n508 7.11588
R3024 vdd.n545 vdd.n536 7.11588
R3025 vdd.n536 vdd.n496 7.11588
R3026 vdd.n668 vdd.n516 7.11588
R3027 vdd.n668 vdd.n496 7.11588
R3028 vdd.n523 vdd.n515 7.11588
R3029 vdd.n523 vdd.n508 7.11588
R3030 vdd.n520 vdd.n519 7.11588
R3031 vdd.n519 vdd.n508 7.11588
R3032 vdd.n567 vdd.n524 7.11588
R3033 vdd.n524 vdd.n496 7.11588
R3034 vdd.n777 vdd.n776 7.11588
R3035 vdd.n776 vdd.n47 7.11588
R3036 vdd.n59 vdd.n58 7.11588
R3037 vdd.n68 vdd.n59 7.11588
R3038 vdd.n67 vdd.n66 7.11588
R3039 vdd.n68 vdd.n67 7.11588
R3040 vdd.n773 vdd.n80 7.11588
R3041 vdd.n80 vdd.n47 7.11588
R3042 vdd.n798 vdd.n12 7.11588
R3043 vdd.n817 vdd.n12 7.11588
R3044 vdd.n804 vdd.n803 7.11588
R3045 vdd.n803 vdd.n29 7.11588
R3046 vdd.n34 vdd.n33 7.11588
R3047 vdd.n33 vdd.n29 7.11588
R3048 vdd.n819 vdd.n818 7.11588
R3049 vdd.n818 vdd.n817 7.11588
R3050 vdd.n657 vdd 6.74008
R3051 vdd.n824 vdd 6.737
R3052 vdd vdd.n657 6.73352
R3053 vdd.n766 vdd.n1 6.63939
R3054 vdd.n652 vdd.n571 6.63939
R3055 vdd.n590 vdd.n586 5.78175
R3056 vdd.n587 vdd.n585 5.78175
R3057 vdd.n585 vdd.n584 5.78175
R3058 vdd.n615 vdd.n603 5.78175
R3059 vdd.n638 vdd.n603 5.78175
R3060 vdd.n629 vdd.n628 5.78175
R3061 vdd.n628 vdd.n606 5.78175
R3062 vdd.n624 vdd.n623 5.78175
R3063 vdd.n624 vdd.n606 5.78175
R3064 vdd.n621 vdd.n580 5.78175
R3065 vdd.n644 vdd.n580 5.78175
R3066 vdd.n643 vdd.n642 5.78175
R3067 vdd.n644 vdd.n643 5.78175
R3068 vdd.n639 vdd.n605 5.78175
R3069 vdd.n639 vdd.n638 5.78175
R3070 vdd.n699 vdd.n483 5.78175
R3071 vdd.n483 vdd.n454 5.78175
R3072 vdd.n704 vdd.n698 5.78175
R3073 vdd.n698 vdd.n462 5.78175
R3074 vdd.n697 vdd.n478 5.78175
R3075 vdd.n697 vdd.n462 5.78175
R3076 vdd.n730 vdd.n729 5.78175
R3077 vdd.n729 vdd.n454 5.78175
R3078 vdd.n479 vdd.n473 5.78175
R3079 vdd.n473 vdd.n464 5.78175
R3080 vdd.n737 vdd.n472 5.78175
R3081 vdd.n472 vdd.n464 5.78175
R3082 vdd.n470 vdd.n458 5.78175
R3083 vdd.n470 vdd.n464 5.78175
R3084 vdd.n693 vdd.n469 5.78175
R3085 vdd.n469 vdd.n464 5.78175
R3086 vdd.n676 vdd.n507 5.78175
R3087 vdd.n676 vdd.n675 5.78175
R3088 vdd.n544 vdd.n505 5.78175
R3089 vdd.n675 vdd.n505 5.78175
R3090 vdd.n719 vdd.n692 5.78175
R3091 vdd.n692 vdd.n454 5.78175
R3092 vdd.n709 vdd.n466 5.78175
R3093 vdd.n709 vdd.n462 5.78175
R3094 vdd.n714 vdd.n713 5.78175
R3095 vdd.n713 vdd.n462 5.78175
R3096 vdd.n716 vdd.n691 5.78175
R3097 vdd.n691 vdd.n454 5.78175
R3098 vdd.n504 vdd.n498 5.78175
R3099 vdd.n683 vdd.n498 5.78175
R3100 vdd.n551 vdd.n542 5.78175
R3101 vdd.n552 vdd.n551 5.78175
R3102 vdd.n554 vdd.n553 5.78175
R3103 vdd.n553 vdd.n552 5.78175
R3104 vdd.n682 vdd.n681 5.78175
R3105 vdd.n683 vdd.n682 5.78175
R3106 vdd.n531 vdd.n497 5.78175
R3107 vdd.n683 vdd.n497 5.78175
R3108 vdd.n527 vdd.n489 5.78175
R3109 vdd.n552 vdd.n489 5.78175
R3110 vdd.n528 vdd.n509 5.78175
R3111 vdd.n675 vdd.n509 5.78175
R3112 vdd.n685 vdd.n684 5.78175
R3113 vdd.n684 vdd.n683 5.78175
R3114 vdd.n687 vdd.n490 5.78175
R3115 vdd.n552 vdd.n490 5.78175
R3116 vdd.n674 vdd.n673 5.78175
R3117 vdd.n675 vdd.n674 5.78175
R3118 vdd.n785 vdd.n40 5.78175
R3119 vdd.n74 vdd.n40 5.78175
R3120 vdd.n57 vdd.n42 5.78175
R3121 vdd.n69 vdd.n57 5.78175
R3122 vdd.n71 vdd.n70 5.78175
R3123 vdd.n70 vdd.n69 5.78175
R3124 vdd.n78 vdd.n39 5.78175
R3125 vdd.n74 vdd.n39 5.78175
R3126 vdd.n73 vdd.n72 5.78175
R3127 vdd.n73 vdd.n46 5.78175
R3128 vdd.n52 vdd.n51 5.78175
R3129 vdd.n52 vdd.n46 5.78175
R3130 vdd.n816 vdd.n815 5.78175
R3131 vdd.n807 vdd.n806 5.78175
R3132 vdd.n808 vdd.n807 5.78175
R3133 vdd.n794 vdd.n18 5.78175
R3134 vdd.n795 vdd.n794 5.78175
R3135 vdd.n24 vdd.n13 5.78175
R3136 vdd.n816 vdd.n13 5.78175
R3137 vdd.n809 vdd.n27 5.78175
R3138 vdd.n809 vdd.n808 5.78175
R3139 vdd.n797 vdd.n796 5.78175
R3140 vdd.n796 vdd.n795 5.78175
R3141 vdd.n21 vdd.n8 4.93648
R3142 vdd.n595 vdd.n590 4.71629
R3143 vdd.n602 vdd.n575 4.7119
R3144 vdd.n679 vdd.n503 4.7119
R3145 vdd.n534 vdd.n533 4.7119
R3146 vdd.n724 vdd.n718 4.7119
R3147 vdd.n484 vdd.n448 4.7119
R3148 vdd.n774 vdd.n41 4.7119
R3149 vdd.n634 vdd.n633 4.70083
R3150 vdd.n557 vdd.n556 4.70083
R3151 vdd.n521 vdd.n491 4.70083
R3152 vdd.n468 vdd.n467 4.70083
R3153 vdd.n477 vdd.n476 4.70083
R3154 vdd.n37 vdd.n36 4.70083
R3155 vdd.n65 vdd.n64 4.70083
R3156 vdd.n588 vdd.n586 4.37746
R3157 vdd.n644 vdd.n581 3.98297
R3158 vdd.n464 vdd.n451 3.98297
R3159 vdd.n675 vdd.n512 3.98297
R3160 vdd.n75 vdd.n74 3.98297
R3161 vdd.n816 vdd.n14 3.98297
R3162 vdd.n569 vdd 3.52106
R3163 vdd.n762 vdd 3.52106
R3164 vdd.n763 vdd.n443 3.32168
R3165 vdd vdd.n168 3.05185
R3166 vdd.n572 vdd 2.62366
R3167 vdd.n398 vdd 2.3405
R3168 vdd.n398 vdd 2.3405
R3169 vdd.n428 vdd 2.3405
R3170 vdd.n428 vdd 2.3405
R3171 vdd.n146 vdd 2.3405
R3172 vdd.n145 vdd 2.3405
R3173 vdd.n104 vdd 2.3405
R3174 vdd.n106 vdd 2.3405
R3175 vdd.n266 vdd 2.3405
R3176 vdd.n266 vdd 2.3405
R3177 vdd.n312 vdd 2.3405
R3178 vdd.n312 vdd 2.3405
R3179 vdd.n214 vdd 2.3405
R3180 vdd.n214 vdd 2.3405
R3181 vdd.n186 vdd 2.3405
R3182 vdd.n186 vdd 2.3405
R3183 vdd.n354 vdd 2.3405
R3184 vdd.n354 vdd 2.3405
R3185 vdd.n384 vdd 2.3405
R3186 vdd.n384 vdd 2.3405
R3187 vdd.n82 vdd 2.29412
R3188 vdd.n313 vdd 2.29412
R3189 vdd.n171 vdd 2.29412
R3190 vdd.n171 vdd 2.29412
R3191 vdd.n721 vdd.n454 1.99173
R3192 vdd.n683 vdd.n499 1.99173
R3193 vdd.n446 vdd 1.93224
R3194 vdd.n660 vdd 1.93224
R3195 vdd.n107 vdd.n106 1.92169
R3196 vdd.n823 vdd 1.89811
R3197 vdd.n767 vdd 1.89811
R3198 vdd.n438 vdd.n397 1.8605
R3199 vdd.n429 vdd.n427 1.8605
R3200 vdd.n438 vdd.n437 1.8605
R3201 vdd.n430 vdd.n429 1.8605
R3202 vdd.n105 vdd.n99 1.8605
R3203 vdd.n144 vdd.n139 1.8605
R3204 vdd.n148 vdd.n147 1.8605
R3205 vdd.n267 vdd.n261 1.8605
R3206 vdd.n311 vdd.n249 1.8605
R3207 vdd.n215 vdd.n184 1.8605
R3208 vdd.n213 vdd.n185 1.8605
R3209 vdd.n268 vdd.n267 1.8605
R3210 vdd.n311 vdd.n310 1.8605
R3211 vdd.n216 vdd.n215 1.8605
R3212 vdd.n213 vdd.n212 1.8605
R3213 vdd.n394 vdd.n353 1.8605
R3214 vdd.n385 vdd.n383 1.8605
R3215 vdd.n394 vdd.n393 1.8605
R3216 vdd.n386 vdd.n385 1.8605
R3217 vdd.n631 vdd.n629 1.77828
R3218 vdd.n559 vdd.n542 1.77828
R3219 vdd.n745 vdd.n466 1.77828
R3220 vdd.n739 vdd.n478 1.77828
R3221 vdd.n527 vdd.n526 1.77828
R3222 vdd.n71 vdd.n54 1.77828
R3223 vdd.n806 vdd.n805 1.77828
R3224 vdd.n351 vdd.n169 1.76063
R3225 vdd.n440 vdd.n439 1.76063
R3226 vdd.n656 vdd.n655 1.753
R3227 vdd.n654 vdd.n570 1.753
R3228 vdd.n396 vdd.n395 1.75125
R3229 vdd.n827 vdd.n826 1.603
R3230 vdd.n825 vdd.n0 1.603
R3231 vdd.n797 vdd.n32 1.5976
R3232 vdd.n650 vdd 1.43984
R3233 vdd.n588 vdd.n584 1.40064
R3234 vdd.n654 vdd.n653 1.35732
R3235 vdd.n617 vdd.n615 1.3042
R3236 vdd.n547 vdd.n544 1.3042
R3237 vdd.n694 vdd.n693 1.3042
R3238 vdd.n480 vdd.n479 1.3042
R3239 vdd.n529 vdd.n528 1.3042
R3240 vdd.n72 vdd.n43 1.3042
R3241 vdd.n813 vdd.n18 1.3042
R3242 vdd.n352 vdd.n351 1.28995
R3243 vdd.n608 vdd.n605 1.19372
R3244 vdd.n539 vdd.n507 1.19372
R3245 vdd.n753 vdd.n458 1.19372
R3246 vdd.n737 vdd.n736 1.19372
R3247 vdd.n673 vdd.n672 1.19372
R3248 vdd.n778 vdd.n51 1.19372
R3249 vdd.n799 vdd.n797 1.19372
R3250 vdd.n395 vdd.n352 1.06531
R3251 vdd.n573 vdd 1.06379
R3252 vdd.n439 vdd.n438 1.06168
R3253 vdd.n395 vdd.n394 1.06168
R3254 vdd.n439 vdd.n81 1.05594
R3255 vdd.n770 vdd 1.04172
R3256 vdd.n6 vdd 1.04172
R3257 vdd.n441 vdd.n81 0.974078
R3258 vdd.n764 vdd.n442 0.918935
R3259 vdd.n761 vdd 0.890303
R3260 vdd.n566 vdd 0.890303
R3261 vdd.n441 vdd.n440 0.855704
R3262 vdd.n591 vdd 0.85529
R3263 vdd.n768 vdd 0.854351
R3264 vdd.n822 vdd 0.854351
R3265 vdd.n765 vdd.n764 0.781762
R3266 vdd.n571 vdd 0.768852
R3267 vdd.n167 vdd.n166 0.715885
R3268 vdd.n349 vdd.n170 0.715885
R3269 vdd.n315 vdd.n314 0.715885
R3270 vdd.n349 vdd.n348 0.715885
R3271 vdd.n824 vdd 0.69425
R3272 vdd.n766 vdd 0.69425
R3273 vdd.n651 vdd.n650 0.619997
R3274 vdd.n573 vdd.n572 0.619997
R3275 vdd.n765 vdd 0.559955
R3276 vdd.n446 vdd.n445 0.518921
R3277 vdd.n762 vdd.n761 0.518921
R3278 vdd.n569 vdd.n566 0.518921
R3279 vdd.n660 vdd.n659 0.518921
R3280 vdd.n443 vdd 0.505434
R3281 vdd.n658 vdd 0.505434
R3282 vdd.n770 vdd.n769 0.497975
R3283 vdd.n768 vdd.n767 0.497975
R3284 vdd.n823 vdd.n822 0.497975
R3285 vdd.n655 vdd.n0 0.479286
R3286 vdd.n763 vdd 0.467672
R3287 vdd.n657 vdd 0.467461
R3288 vdd.n168 vdd 0.464224
R3289 vdd.n764 vdd.n763 0.426664
R3290 vdd.n314 vdd 0.413
R3291 vdd.n350 vdd.n349 0.410656
R3292 vdd.n648 vdd.n574 0.376971
R3293 vdd.n431 vdd.n430 0.376971
R3294 vdd.n437 vdd.n399 0.376971
R3295 vdd.n427 vdd.n410 0.376971
R3296 vdd.n420 vdd.n397 0.376971
R3297 vdd.n148 vdd.n143 0.376971
R3298 vdd.n139 vdd.n138 0.376971
R3299 vdd.n166 vdd.n83 0.376971
R3300 vdd.n100 vdd.n99 0.376971
R3301 vdd.n108 vdd.n107 0.376971
R3302 vdd.n662 vdd.n565 0.376971
R3303 vdd.n459 vdd.n444 0.376971
R3304 vdd.n759 vdd.n447 0.376971
R3305 vdd.n568 vdd.n517 0.376971
R3306 vdd.n772 vdd.n50 0.376971
R3307 vdd.n820 vdd.n7 0.376971
R3308 vdd.n212 vdd.n187 0.376971
R3309 vdd.n217 vdd.n216 0.376971
R3310 vdd.n348 vdd.n172 0.376971
R3311 vdd.n315 vdd.n248 0.376971
R3312 vdd.n310 vdd.n250 0.376971
R3313 vdd.n269 vdd.n268 0.376971
R3314 vdd.n193 vdd.n185 0.376971
R3315 vdd.n196 vdd.n184 0.376971
R3316 vdd.n338 vdd.n170 0.376971
R3317 vdd.n256 vdd.n249 0.376971
R3318 vdd.n262 vdd.n261 0.376971
R3319 vdd.n387 vdd.n386 0.376971
R3320 vdd.n393 vdd.n355 0.376971
R3321 vdd.n383 vdd.n366 0.376971
R3322 vdd.n376 vdd.n353 0.376971
R3323 vdd.n652 vdd 0.376726
R3324 vdd.n314 vdd.n313 0.360656
R3325 vdd.n349 vdd.n171 0.360656
R3326 vdd.n591 vdd 0.349949
R3327 vdd.n593 vdd 0.344944
R3328 vdd.n442 vdd.n441 0.34097
R3329 vdd.n632 vdd.n631 0.307571
R3330 vdd.n559 vdd.n558 0.307571
R3331 vdd.n745 vdd.n744 0.307571
R3332 vdd.n740 vdd.n739 0.307571
R3333 vdd.n526 vdd.n525 0.307571
R3334 vdd.n63 vdd.n54 0.307571
R3335 vdd.n805 vdd.n30 0.307571
R3336 vdd.n651 vdd 0.304352
R3337 vdd.n595 vdd.n594 0.291125
R3338 vdd.n593 vdd.n592 0.277007
R3339 vdd.n1 vdd 0.27355
R3340 vdd.n594 vdd.n591 0.2731
R3341 vdd.n2 vdd 0.272663
R3342 vdd.n440 vdd.n396 0.264604
R3343 vdd.n396 vdd.n169 0.263158
R3344 vdd.n445 vdd 0.254776
R3345 vdd.n659 vdd 0.254776
R3346 vdd.n6 vdd.n5 0.249237
R3347 vdd.n5 vdd.n3 0.249237
R3348 vdd.n769 vdd 0.244503
R3349 vdd.n3 vdd 0.244503
R3350 vdd.n352 vdd.n81 0.233429
R3351 vdd.n168 vdd.n167 0.22821
R3352 vdd.n167 vdd.n82 0.201986
R3353 vdd.n642 vdd.n641 0.178728
R3354 vdd.n678 vdd.n504 0.178728
R3355 vdd.n723 vdd.n719 0.178728
R3356 vdd.n730 vdd.n481 0.178728
R3357 vdd.n532 vdd.n531 0.178728
R3358 vdd.n78 vdd.n77 0.178728
R3359 vdd.n215 vdd 0.166125
R3360 vdd.n429 vdd 0.164562
R3361 vdd.n311 vdd 0.164562
R3362 vdd vdd.n213 0.164562
R3363 vdd.n385 vdd 0.164562
R3364 vdd vdd.n824 0.148
R3365 vdd.n761 vdd.n760 0.147704
R3366 vdd.n661 vdd.n566 0.147704
R3367 vdd.n760 vdd.n446 0.146059
R3368 vdd.n661 vdd.n660 0.146059
R3369 vdd.n649 vdd.n648 0.133357
R3370 vdd.n760 vdd.n444 0.133357
R3371 vdd.n760 vdd.n759 0.133357
R3372 vdd.n661 vdd.n568 0.133357
R3373 vdd.n662 vdd.n661 0.133357
R3374 vdd.n772 vdd.n771 0.133357
R3375 vdd.n821 vdd.n820 0.133357
R3376 vdd.n445 vdd.n443 0.131257
R3377 vdd.n659 vdd.n658 0.131257
R3378 vdd.n763 vdd.n762 0.131257
R3379 vdd.n657 vdd.n569 0.129612
R3380 vdd.n592 vdd 0.113524
R3381 vdd.n649 vdd.n573 0.110181
R3382 vdd.n438 vdd.n398 0.109875
R3383 vdd.n429 vdd.n428 0.109875
R3384 vdd.n267 vdd.n266 0.109875
R3385 vdd.n312 vdd.n311 0.109875
R3386 vdd.n215 vdd.n214 0.109875
R3387 vdd.n213 vdd.n186 0.109875
R3388 vdd.n394 vdd.n354 0.109875
R3389 vdd.n385 vdd.n384 0.109875
R3390 vdd.n650 vdd.n649 0.108956
R3391 vdd.n657 vdd 0.100037
R3392 vdd.n652 vdd.n651 0.0979265
R3393 vdd.n642 vdd.n601 0.0977152
R3394 vdd.n546 vdd.n504 0.0977152
R3395 vdd.n719 vdd.n457 0.0977152
R3396 vdd.n731 vdd.n730 0.0977152
R3397 vdd.n531 vdd.n530 0.0977152
R3398 vdd.n79 vdd.n78 0.0977152
R3399 vdd.n572 vdd.n571 0.096701
R3400 vdd.n144 vdd 0.0931573
R3401 vdd vdd.n105 0.0922832
R3402 vdd.n147 vdd 0.0922832
R3403 vdd.n592 vdd 0.0847634
R3404 vdd.n771 vdd.n768 0.079844
R3405 vdd.n822 vdd.n821 0.079844
R3406 vdd.n771 vdd.n770 0.0789574
R3407 vdd.n821 vdd.n6 0.0789574
R3408 vdd.n351 vdd.n350 0.0780862
R3409 vdd.n3 vdd.n2 0.0709787
R3410 vdd.n824 vdd.n823 0.0709787
R3411 vdd.n767 vdd.n766 0.0709787
R3412 vdd.n769 vdd.n1 0.0700922
R3413 vdd.n653 vdd 0.0630773
R3414 vdd.n105 vdd.n104 0.0616888
R3415 vdd.n145 vdd.n144 0.0616888
R3416 vdd.n147 vdd.n146 0.0616888
R3417 vdd.n571 vdd.n442 0.0572867
R3418 vdd vdd.n398 0.0551875
R3419 vdd.n428 vdd 0.0551875
R3420 vdd.n266 vdd 0.0551875
R3421 vdd vdd.n312 0.0551875
R3422 vdd.n214 vdd 0.0551875
R3423 vdd.n186 vdd 0.0551875
R3424 vdd vdd.n354 0.0551875
R3425 vdd.n384 vdd 0.0551875
R3426 vdd.n825 vdd 0.0545625
R3427 vdd.n313 vdd 0.0512812
R3428 vdd vdd.n171 0.0512812
R3429 vdd.n653 vdd.n652 0.045162
R3430 vdd.n655 vdd.n654 0.0388531
R3431 vdd.n826 vdd.n1 0.0351875
R3432 vdd vdd.n656 0.0334335
R3433 vdd.n570 vdd.n443 0.0315396
R3434 vdd.n106 vdd 0.0310944
R3435 vdd.n104 vdd 0.0310944
R3436 vdd vdd.n145 0.0310944
R3437 vdd.n146 vdd 0.0310944
R3438 vdd.n766 vdd.n765 0.0298951
R3439 vdd vdd.n82 0.0289091
R3440 vdd.n2 vdd 0.0265417
R3441 vdd.n827 vdd.n0 0.0256039
R3442 vdd.n658 vdd 0.0140031
R3443 vdd.n826 vdd.n825 0.008
R3444 vdd.n658 vdd 0.00744444
R3445 vdd.n169 vdd 0.00538077
R3446 vdd.n594 vdd.n593 0.00440625
R3447 vdd vdd.n827 0.00308012
R3448 vdd.n350 vdd 0.00284375
R3449 vdd.n656 vdd.n570 0.00113131
R3450 vref.n0 vref 2.51601
R3451 vref.n0 vref 2.11902
R3452 vref vref.n1 1.37411
R3453 vref.n1 vref 0.831056
R3454 vref.n1 vref 0.774111
R3455 vref.n1 vref 0.231056
R3456 vref vref.n0 0.188289
R3457 vref.n1 vref 0.0135208
R3458 vref.n1 vref 0.0135208
R3459 comp_p_1/latch_left.n0 comp_p_1/latch_left.t3 114.778
R3460 comp_p_1/latch_left.n0 comp_p_1/latch_left.t2 106.572
R3461 comp_p_1/latch_left.n1 comp_p_1/latch_left.t0 95.1712
R3462 comp_p_1/latch_left.n2 comp_p_1/latch_left.t1 22.0141
R3463 comp_p_1/latch_left.n1 comp_p_1/latch_left.n0 1.72733
R3464 comp_p_1/latch_left comp_p_1/latch_left.n2 0.717514
R3465 comp_p_1/latch_left.n2 comp_p_1/latch_left.n1 0.599169
R3466 d0.n0 d0.t1 556.78
R3467 d0.t1 d0 547.24
R3468 d0 d0.t0 372.113
R3469 d0.n0 d0 9.54008
R3470 d0.n2 d0 6.80006
R3471 d0 d0.n2 4.54809
R3472 d0.n3 d0 0.719145
R3473 d0.n1 d0.n0 0.253625
R3474 d0 d0.n3 0.199411
R3475 d0 d0 0.063
R3476 d0.n2 d0 0.0443144
R3477 d0.n3 d0 0.0262742
R3478 d0 d0 0.0262732
R3479 d0.n1 d0 0.013
R3480 d0.n3 d0 0.00763393
R3481 d0 d0.n1 0.00565464
R3482 vin.n20 vin.t26 899.324
R3483 vin.n38 vin.t22 899.324
R3484 vin.n31 vin.t14 899.324
R3485 vin.n25 vin.t2 899.324
R3486 vin.n2 vin.t6 899.324
R3487 vin.n7 vin.t10 899.324
R3488 vin.n13 vin.t18 899.324
R3489 vin.n21 vin.t26 898.659
R3490 vin.n39 vin.t22 898.659
R3491 vin.n32 vin.t14 898.659
R3492 vin.n26 vin.t2 898.659
R3493 vin.n3 vin.t6 898.659
R3494 vin.n8 vin.t10 898.659
R3495 vin.n14 vin.t18 898.659
R3496 vin.t23 vin.n38 898.442
R3497 vin.t3 vin.n25 898.442
R3498 vin.t7 vin.n2 898.442
R3499 vin.t19 vin.n13 898.442
R3500 vin.t27 vin.n20 898.442
R3501 vin.t15 vin.n31 898.442
R3502 vin.t11 vin.n7 898.442
R3503 vin.n21 vin.t27 897.754
R3504 vin.n39 vin.t23 897.754
R3505 vin.n32 vin.t15 897.754
R3506 vin.n26 vin.t3 897.754
R3507 vin.n3 vin.t7 897.754
R3508 vin.n8 vin.t11 897.754
R3509 vin.n14 vin.t19 897.754
R3510 vin.n18 vin.t24 895.625
R3511 vin.n36 vin.t20 895.625
R3512 vin.n29 vin.t12 895.625
R3513 vin.n23 vin.t0 895.625
R3514 vin.n0 vin.t4 895.625
R3515 vin.n5 vin.t8 895.625
R3516 vin.n11 vin.t16 895.625
R3517 vin.n18 vin.t25 894.172
R3518 vin.n36 vin.t21 894.172
R3519 vin.n29 vin.t13 894.172
R3520 vin.n23 vin.t1 894.172
R3521 vin.n0 vin.t5 894.172
R3522 vin.n5 vin.t9 894.172
R3523 vin.n11 vin.t17 894.172
R3524 vin.n19 vin.n18 6.30807
R3525 vin.n37 vin.n36 6.30807
R3526 vin.n30 vin.n29 6.30807
R3527 vin.n24 vin.n23 6.30807
R3528 vin.n1 vin.n0 6.30807
R3529 vin.n6 vin.n5 6.30807
R3530 vin.n12 vin.n11 6.30807
R3531 vin.n20 vin.n19 5.39021
R3532 vin.n38 vin.n37 5.39021
R3533 vin.n31 vin.n30 5.39021
R3534 vin.n25 vin.n24 5.39021
R3535 vin.n2 vin.n1 5.39021
R3536 vin.n7 vin.n6 5.39021
R3537 vin.n13 vin.n12 5.39021
R3538 vin.n22 vin.n21 5.38653
R3539 vin.n40 vin.n39 5.38653
R3540 vin.n33 vin.n32 5.38653
R3541 vin.n27 vin.n26 5.38653
R3542 vin.n4 vin.n3 5.38653
R3543 vin.n9 vin.n8 5.38653
R3544 vin.n15 vin.n14 5.38653
R3545 vin.n44 vin.n43 5.20469
R3546 vin.n22 vin.n19 5.11108
R3547 vin.n40 vin.n37 5.11108
R3548 vin.n33 vin.n30 5.11108
R3549 vin.n27 vin.n24 5.11108
R3550 vin.n4 vin.n1 5.11108
R3551 vin.n9 vin.n6 5.11108
R3552 vin.n15 vin.n12 5.11108
R3553 vin.n35 vin.n28 4.57467
R3554 vin.n10 vin 4.13219
R3555 vin.n35 vin.n34 3.68222
R3556 vin.n42 vin.n41 3.10272
R3557 vin.n16 vin 2.68025
R3558 vin.n10 vin 2.66582
R3559 vin.n43 vin.n42 2.43775
R3560 vin.n43 vin 1.54614
R3561 vin vin.n16 1.12357
R3562 vin vin.n22 0.870692
R3563 vin vin.n4 0.870692
R3564 vin vin.n9 0.870692
R3565 vin vin.n15 0.870692
R3566 vin.n34 vin.n33 0.837038
R3567 vin.n41 vin.n40 0.726462
R3568 vin.n16 vin.n10 0.70492
R3569 vin.n28 vin.n27 0.668769
R3570 vin.n42 vin.n35 0.533734
R3571 vin.n17 vin 0.468179
R3572 vin vin.n45 0.371278
R3573 vin.n45 vin 0.332981
R3574 vin.n17 vin 0.23608
R3575 vin.n45 vin 0.20608
R3576 vin.n17 vin 0.146164
R3577 vin.n41 vin 0.0482941
R3578 vin.n44 vin.n17 0.0422977
R3579 vin.n45 vin.n44 0.0422977
R3580 vin.n28 vin 0.0391905
R3581 vin.n34 vin 0.0341538
R3582 comp_p_0/latch_right.n1 comp_p_0/latch_right.t3 114.778
R3583 comp_p_0/latch_right.n1 comp_p_0/latch_right.t2 106.572
R3584 comp_p_0/latch_right.n2 comp_p_0/latch_right.t0 94.6192
R3585 comp_p_0/latch_right.n0 comp_p_0/latch_right.t1 22.0141
R3586 comp_p_0/latch_right.n2 comp_p_0/latch_right.n0 2.37533
R3587 comp_p_0/latch_right.n3 comp_p_0/latch_right.n1 1.43373
R3588 comp_p_0/latch_right.n4 comp_p_0/latch_right.n3 1.11841
R3589 comp_p_0/latch_right.n3 comp_p_0/latch_right.n2 1.06963
R3590 comp_p_0/latch_right comp_p_0/latch_right.n4 0.608139
R3591 comp_p_0/latch_right.n4 comp_p_0/latch_right.n0 0.00530769
R3592 comp_p_0/out_left.n1 comp_p_0/out_left.t2 145.612
R3593 comp_p_0/out_left.n2 comp_p_0/out_left.t0 143.417
R3594 comp_p_0/out_left.n0 comp_p_0/out_left.t1 29.4286
R3595 comp_p_0/out_left comp_p_0/out_left.n3 11.6041
R3596 comp_p_0/out_left.n3 comp_p_0/out_left.n2 4.33076
R3597 comp_p_0/out_left.n1 comp_p_0/out_left.n0 2.12634
R3598 comp_p_0/out_left.n2 comp_p_0/out_left.n1 2.04428
R3599 comp_p_0/out_left.n3 comp_p_0/out_left.n0 0.00290385
R3600 d1.n0 d1.t1 556.78
R3601 d1.t1 d1 547.24
R3602 d1 d1.t0 372.113
R3603 d1.n1 d1 20.4858
R3604 d1.n0 d1 9.54008
R3605 d1.n1 d1 4.95991
R3606 d1 d1.n1 3.5178
R3607 d1.n2 d1 1.7016
R3608 d1 d1.n2 0.538602
R3609 d1 d1.n0 0.266125
R3610 d1 d1 0.063
R3611 d1.n2 d1 0.0217258
R3612 d1.n2 d1 0.00721429
R3613 comp_p_2/latch_left.n0 comp_p_2/latch_left.t3 114.778
R3614 comp_p_2/latch_left.n0 comp_p_2/latch_left.t2 106.572
R3615 comp_p_2/latch_left.n1 comp_p_2/latch_left.t0 95.1712
R3616 comp_p_2/latch_left.n2 comp_p_2/latch_left.t1 22.0141
R3617 comp_p_2/latch_left.n1 comp_p_2/latch_left.n0 1.72733
R3618 comp_p_2/latch_left comp_p_2/latch_left.n2 0.717514
R3619 comp_p_2/latch_left.n2 comp_p_2/latch_left.n1 0.599169
R3620 comp_p_2/out_left.n1 comp_p_2/out_left.t2 145.612
R3621 comp_p_2/out_left.n2 comp_p_2/out_left.t0 143.417
R3622 comp_p_2/out_left.n0 comp_p_2/out_left.t1 29.4286
R3623 comp_p_2/out_left comp_p_2/out_left.n3 11.6041
R3624 comp_p_2/out_left.n3 comp_p_2/out_left.n2 4.33076
R3625 comp_p_2/out_left.n1 comp_p_2/out_left.n0 2.12634
R3626 comp_p_2/out_left.n2 comp_p_2/out_left.n1 2.04428
R3627 comp_p_2/out_left.n3 comp_p_2/out_left.n0 0.00290385
R3628 d2.n0 d2.t1 556.78
R3629 d2.t1 d2 547.24
R3630 d2 d2.t0 372.113
R3631 d2.n2 d2 18.5303
R3632 d2.n0 d2 9.54008
R3633 d2.n4 d2 2.94937
R3634 d2.n2 d2 1.06045
R3635 d2.n3 d2.n2 0.853
R3636 d2 d2.n4 0.464536
R3637 d2.n1 d2.n0 0.25675
R3638 d2.n4 d2 0.0929839
R3639 d2 d2 0.063
R3640 d2 d2 0.0329675
R3641 d2.n1 d2 0.009875
R3642 d2.n4 d2.n3 0.00777665
R3643 d2.n3 d2 0.00777665
R3644 d2 d2.n1 0.00537013
R3645 comp_p_3/latch_left.n0 comp_p_3/latch_left.t3 114.778
R3646 comp_p_3/latch_left.n0 comp_p_3/latch_left.t2 106.572
R3647 comp_p_3/latch_left.n1 comp_p_3/latch_left.t0 95.1712
R3648 comp_p_3/latch_left.n2 comp_p_3/latch_left.t1 22.0141
R3649 comp_p_3/latch_left.n1 comp_p_3/latch_left.n0 1.72733
R3650 comp_p_3/latch_left comp_p_3/latch_left.n2 0.717514
R3651 comp_p_3/latch_left.n2 comp_p_3/latch_left.n1 0.599169
R3652 d3.n0 d3.t1 556.78
R3653 d3.t1 d3 547.24
R3654 d3 d3.t0 372.113
R3655 d3.n1 d3 10.0074
R3656 d3.n0 d3 9.54008
R3657 d3.n3 d3 3.8636
R3658 d3.n2 d3.n1 1.978
R3659 d3 d3.n3 1.07938
R3660 d3.n1 d3 0.589103
R3661 d3 d3.n0 0.266125
R3662 d3.n3 d3 0.0975323
R3663 d3 d3 0.063
R3664 d3.n3 d3.n2 0.0223063
R3665 d3.n2 d3 0.00579279
R3666 comp_p_4/out_left.n1 comp_p_4/out_left.t2 145.612
R3667 comp_p_4/out_left.n2 comp_p_4/out_left.t0 143.417
R3668 comp_p_4/out_left.n0 comp_p_4/out_left.t1 29.4286
R3669 comp_p_4/out_left comp_p_4/out_left.n3 11.6041
R3670 comp_p_4/out_left.n3 comp_p_4/out_left.n2 4.33076
R3671 comp_p_4/out_left.n1 comp_p_4/out_left.n0 2.12634
R3672 comp_p_4/out_left.n2 comp_p_4/out_left.n1 2.04428
R3673 comp_p_4/out_left.n3 comp_p_4/out_left.n0 0.00290385
R3674 d4.n0 d4.t1 556.78
R3675 d4.t1 d4 547.24
R3676 d4 d4.t0 372.113
R3677 d4.n1 d4 24.0965
R3678 d4.n0 d4 9.54008
R3679 d4.n2 d4 5.15685
R3680 d4.n1 d4 1.81119
R3681 d4 d4.n1 1.16374
R3682 d4 d4.n2 1.15048
R3683 d4 d4.n0 0.266125
R3684 d4 d4 0.063
R3685 d4.n2 d4 0.00656452
R3686 d4.n2 d4 0.00185252
R3687 comp_p_5/latch_left.n0 comp_p_5/latch_left.t3 114.778
R3688 comp_p_5/latch_left.n0 comp_p_5/latch_left.t2 106.572
R3689 comp_p_5/latch_left.n1 comp_p_5/latch_left.t0 95.1712
R3690 comp_p_5/latch_left.n2 comp_p_5/latch_left.t1 22.0141
R3691 comp_p_5/latch_left.n1 comp_p_5/latch_left.n0 1.72733
R3692 comp_p_5/latch_left comp_p_5/latch_left.n2 0.717514
R3693 comp_p_5/latch_left.n2 comp_p_5/latch_left.n1 0.599169
R3694 comp_p_5/latch_right.n1 comp_p_5/latch_right.t3 114.778
R3695 comp_p_5/latch_right.n1 comp_p_5/latch_right.t2 106.572
R3696 comp_p_5/latch_right.n2 comp_p_5/latch_right.t0 94.6192
R3697 comp_p_5/latch_right.n0 comp_p_5/latch_right.t1 22.0141
R3698 comp_p_5/latch_right.n2 comp_p_5/latch_right.n0 2.37533
R3699 comp_p_5/latch_right.n3 comp_p_5/latch_right.n1 1.43373
R3700 comp_p_5/latch_right.n4 comp_p_5/latch_right.n3 1.11841
R3701 comp_p_5/latch_right.n3 comp_p_5/latch_right.n2 1.06963
R3702 comp_p_5/latch_right comp_p_5/latch_right.n4 0.608139
R3703 comp_p_5/latch_right.n4 comp_p_5/latch_right.n0 0.00530769
R3704 d5.n0 d5.t1 556.78
R3705 d5.t1 d5 547.24
R3706 d5 d5.t0 372.113
R3707 d5.n0 d5 9.54008
R3708 d5.n2 d5.n1 7.93228
R3709 d5.n1 d5 7.34675
R3710 d5.n3 d5 6.13627
R3711 d5 d5.n3 1.18931
R3712 d5.n1 d5 0.520292
R3713 d5 d5.n0 0.266125
R3714 d5 d5 0.063
R3715 d5.n3 d5 0.0535645
R3716 d5.n3 d5.n2 0.00564062
R3717 d5.n2 d5 0.00564062
R3718 comp_p_6/out_left.n1 comp_p_6/out_left.t2 145.612
R3719 comp_p_6/out_left.n2 comp_p_6/out_left.t0 143.417
R3720 comp_p_6/out_left.n0 comp_p_6/out_left.t1 29.4286
R3721 comp_p_6/out_left comp_p_6/out_left.n3 11.6041
R3722 comp_p_6/out_left.n3 comp_p_6/out_left.n2 4.33076
R3723 comp_p_6/out_left.n1 comp_p_6/out_left.n0 2.12634
R3724 comp_p_6/out_left.n2 comp_p_6/out_left.n1 2.04428
R3725 comp_p_6/out_left.n3 comp_p_6/out_left.n0 0.00290385
R3726 d6.n0 d6.t1 556.78
R3727 d6.t1 d6 547.24
R3728 d6 d6.t0 372.113
R3729 d6.n1 d6 11.4942
R3730 d6.n0 d6 9.54008
R3731 d6 d6.n2 7.42498
R3732 d6.n2 d6.n1 3.89032
R3733 d6.n1 d6 1.33473
R3734 d6 d6.n0 0.266125
R3735 d6 d6 0.063
R3736 d6.n2 d6 0.0232419
R3737 dout0 dout0 5.30089
R3738 dout0 dout0 2.61734
R3739 dout1 dout1 5.30089
R3740 dout1 dout1 2.61734
R3741 dout2 dout2 5.30089
R3742 dout2 dout2 2.61734
C0 comp_p_0/out_left vin 0.0787f
C1 comp_p_4/latch_left comp_p_4/vinn 0.00288f
C2 d4 comp_p_6/latch_right 0.06065f
C3 d5 d2 0.04522f
C4 comp_p_1/vinn d4 0
C5 comp_p_1/vinn d1 0.26283f
C6 comp_p_1/latch_right d6 0.00271f
C7 vdd comp_p_1/tail 0.35563f
C8 comp_p_1/latch_left comp_p_3/latch_left 0.00925f
C9 comp_p_1/vinn comp_p_6/vbias_p 0.38594f
C10 vin vref 0.01522f
C11 comp_p_0/latch_left comp_p_2/latch_left 0.01494f
C12 vin comp_p_3/out_left 0.05071f
C13 comp_p_6/latch_left vbias_generation_0/bias_n 0.01259f
C14 vin vdd 10.42758f
C15 d4 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00277f
C16 d5 d4 4.7254f
C17 d5 d1 0.06814f
C18 d5 comp_p_6/vbias_p 0.00462f
C19 comp_p_4/latch_right vdd 0.00589f
C20 vin comp_p_0/vinn 0.81463f
C21 comp_p_6/tail vdd 0.35623f
C22 comp_p_2/latch_right comp_p_3/out_left 0
C23 comp_p_2/latch_right vdd 0.00592f
C24 vin vbias_generation_0/XR_bias_3/R2 0.08368f
C25 comp_p_1/vinn d3 0
C26 comp_p_6/vinn vbias_generation_0/bias_n 0.43753f
C27 comp_p_6/tail vbias_generation_0/XR_bias_3/R2 0
C28 d5 comp_p_3/tail 0
C29 d5 d3 0.16529f
C30 comp_p_4/vinn comp_p_5/out_left 0
C31 d2 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C32 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G d0 0
C33 tmux_7therm_to_3bin_0/buffer_4/out vdd 0.00843f
C34 comp_p_1/vinn vin 0.95805f
C35 comp_p_5/vinn comp_p_3/vinn 0.0226f
C36 d4 tmux_7therm_to_3bin_0/buffer_5/out 0.01207f
C37 comp_p_3/out_left comp_p_2/vinn 0
C38 d5 comp_p_1/tail 0
C39 comp_p_2/vinn vdd 0.04727f
C40 d4 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0.00187f
C41 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vdd 0.00104f
C42 d4 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C43 d1 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0.00131f
C44 d5 vin 0.0056f
C45 comp_p_6/out_left vdd 1.84652f
C46 comp_p_1/vinn comp_p_2/latch_right 0.00771f
C47 comp_p_1/out_left d6 0
C48 comp_p_6/vbias_p comp_p_4/out_left 0.69034f
C49 comp_p_2/vinn comp_p_0/vinn 0.02754f
C50 comp_p_5/latch_left comp_p_6/latch_left 0.00925f
C51 comp_p_1/latch_right vdd 1.96641f
C52 d0 d6 0.07778f
C53 vbias_generation_0/XR_bias_4/R1 comp_p_6/vinn 0.51064f
C54 comp_p_6/out_left vbias_generation_0/XR_bias_3/R2 0.00563f
C55 d4 comp_p_5/vinn 0.25745f
C56 comp_p_6/vinn comp_p_6/latch_left 0.00473f
C57 comp_p_6/vbias_p comp_p_5/vinn 0.407f
C58 d3 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C59 d5 tmux_7therm_to_3bin_0/buffer_4/out 0
C60 comp_p_0/latch_right vdd 0.00588f
C61 tmux_7therm_to_3bin_0/R1/R1 vdd 0.00399f
C62 d2 tmux_7therm_to_3bin_0/buffer_0/out 0
C63 tmux_7therm_to_3bin_0/tmux_2to1_3/A d0 0
C64 vin comp_p_4/out_left 0.0859f
C65 d5 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin 0
C66 comp_p_1/vinn comp_p_1/latch_right 0.00799f
C67 comp_p_0/latch_right comp_p_0/vinn 0.00236f
C68 comp_p_5/latch_left d6 0.00183f
C69 comp_p_6/vbias_p comp_p_4/latch_left 0.37827f
C70 comp_p_0/latch_left vdd 0
C71 d4 tmux_7therm_to_3bin_0/buffer_0/out 0
C72 d1 tmux_7therm_to_3bin_0/buffer_0/out 0
C73 vdd vbias_generation_0/bias_n 0.0189f
C74 d5 comp_p_1/latch_right 0.0019f
C75 vin comp_p_5/vinn 0.66275f
C76 comp_p_0/latch_left comp_p_0/vinn 0.02494f
C77 comp_p_1/latch_left d2 0
C78 comp_p_5/latch_right d6 0
C79 comp_p_1/out_left vdd 1.79183f
C80 comp_p_4/latch_right comp_p_5/vinn 0.20935f
C81 comp_p_3/vinn comp_p_3/latch_left 0.00666f
C82 comp_p_1/vinn comp_p_0/latch_right 0.1958f
C83 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d2 0.00484f
C84 d4 comp_p_1/latch_left 0
C85 comp_p_1/latch_left d1 0.09499f
C86 d0 vdd 2.70776f
C87 comp_p_1/out_left comp_p_0/vinn 0
C88 tmux_7therm_to_3bin_0/buffer_0/out d3 0
C89 comp_p_3/vinn comp_p_3/latch_right 0.00805f
C90 vbias_generation_0/XR_bias_2/R2 comp_p_6/vbias_p 0.02749f
C91 d2 comp_p_3/latch_left 0.09614f
C92 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin d6 0
C93 d4 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C94 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d1 0.00256f
C95 comp_p_0/latch_left comp_p_1/vinn 0.15776f
C96 d4 comp_p_5/out_left 0.61143f
C97 vin comp_p_4/latch_left 0.00664f
C98 comp_p_6/vbias_p comp_p_5/out_left -0.0642f
C99 comp_p_6/latch_right vbias_generation_0/bias_n 0
C100 d2 comp_p_3/latch_right 0.09517f
C101 comp_p_3/vinn comp_p_4/vinn 0
C102 d1 comp_p_3/latch_left 0
C103 d4 comp_p_3/latch_left 0
C104 comp_p_0/out_left comp_p_2/latch_left 0.01472f
C105 comp_p_3/vinn comp_p_2/out_left 0.01462f
C106 d4 comp_p_5/tail 0.00266f
C107 comp_p_1/latch_left d3 0
C108 comp_p_1/vinn comp_p_1/out_left 0.19389f
C109 vdd comp_p_4/tail 0.00166f
C110 d1 comp_p_3/latch_right 0
C111 d4 comp_p_3/latch_right 0.00133f
C112 comp_p_6/latch_left vdd 2.00132f
C113 comp_p_2/latch_left vdd 0
C114 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d3 0
C115 comp_p_5/latch_left vdd 2.04609f
C116 d3 comp_p_5/out_left 0.02309f
C117 d5 comp_p_1/out_left 0
C118 vdd tmux_7therm_to_3bin_0/buffer_8/in 0
C119 d4 comp_p_4/vinn -0
C120 comp_p_2/latch_left comp_p_0/vinn 0
C121 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vdd 0.00166f
C122 comp_p_6/vinn vref 0.00148f
C123 comp_p_6/vbias_p comp_p_4/vinn 0.12306f
C124 d3 comp_p_3/latch_left 0
C125 vbias_generation_0/XR_bias_2/R2 vin 0.50675f
C126 d5 d0 0.04624f
C127 comp_p_6/vinn vdd 1.11418f
C128 comp_p_6/vbias_p comp_p_2/out_left 0.68901f
C129 comp_p_5/latch_right vdd 1.9557f
C130 d3 comp_p_3/latch_right 0.0057f
C131 vin comp_p_5/out_left 0.06043f
C132 comp_p_4/latch_right comp_p_5/out_left 0
C133 d2 tmux_7therm_to_3bin_0/buffer_1/out 0
C134 comp_p_6/vinn vbias_generation_0/XR_bias_3/R2 0.06411f
C135 vin comp_p_5/tail 0.00233f
C136 comp_p_3/out_left d6 0
C137 comp_p_1/vinn comp_p_2/latch_left 0.01672f
C138 comp_p_2/tail comp_p_3/out_left 0
C139 comp_p_0/tail d1 -0.00224f
C140 vdd d6 5.14584f
C141 comp_p_2/tail vdd 0.00168f
C142 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin vdd 0
C143 comp_p_0/tail comp_p_6/vbias_p 0.31444f
C144 d2 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0.00171f
C145 d1 tmux_7therm_to_3bin_0/buffer_1/out 0.01519f
C146 comp_p_2/latch_right comp_p_3/latch_left 0.02598f
C147 comp_p_6/vinn comp_p_6/latch_right 0.00296f
C148 vin comp_p_4/vinn 0.52728f
C149 d4 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C150 d1 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0.00562f
C151 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d0 0.00746f
C152 comp_p_5/latch_right comp_p_6/latch_right 0.00925f
C153 vin comp_p_2/out_left 0.0842f
C154 d3 tmux_7therm_to_3bin_0/R1/R2 0
C155 comp_p_4/latch_right comp_p_4/vinn 0.00144f
C156 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vdd 0.00166f
C157 tmux_7therm_to_3bin_0/tmux_2to1_3/A vdd 0.00153f
C158 comp_p_1/vinn d6 0
C159 comp_p_3/vinn d2 0.24742f
C160 vbias_generation_0/XR_bias_4/R1 comp_p_4/out_left 0
C161 d3 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C162 comp_p_0/tail vin 0.01181f
C163 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin d6 0
C164 comp_p_4/latch_left vbias_generation_0/bias_n 0
C165 d5 d6 4.41099f
C166 d5 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C167 d4 comp_p_3/vinn 0
C168 comp_p_0/out_left vdd 0.01217f
C169 comp_p_3/vinn d1 0
C170 comp_p_6/vbias_p comp_p_3/vinn 0.38072f
C171 comp_p_0/latch_right comp_p_1/latch_left 0.02598f
C172 d4 tmux_7therm_to_3bin_0/buffer_6/out 0.01165f
C173 comp_p_1/latch_right comp_p_3/latch_right 0.00925f
C174 comp_p_0/out_left comp_p_0/vinn 0.02276f
C175 comp_p_3/out_left vdd 1.79594f
C176 comp_p_2/out_left comp_p_2/vinn 0.0232f
C177 d4 d2 0.0466f
C178 comp_p_5/vinn comp_p_4/tail 0.10856f
C179 d2 d1 3.65092f
C180 d1 tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G 0
C181 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin tmux_7therm_to_3bin_0/R1/R1 -0
C182 comp_p_6/vbias_p d2 0.37534f
C183 comp_p_6/vinn comp_p_4/out_left 0.04948f
C184 tmux_7therm_to_3bin_0/buffer_0/out d0 0
C185 comp_p_5/latch_left comp_p_5/vinn 0.00674f
C186 vdd comp_p_0/vinn 0.01961f
C187 comp_p_3/vinn d3 0.0076f
C188 d4 d1 0.10688f
C189 vbias_generation_0/XR_bias_3/R2 vdd 0.08059f
C190 d4 comp_p_6/vbias_p 0.37293f
C191 comp_p_6/vbias_p d1 0.37529f
C192 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin d6 0.00531f
C193 comp_p_1/vinn comp_p_0/out_left 0.03983f
C194 comp_p_6/vinn comp_p_5/vinn 0.03037f
C195 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin d6 0
C196 vbias_generation_0/XR_bias_4/R1 comp_p_4/latch_left 0
C197 comp_p_3/tail d2 0.00272f
C198 d2 d3 2.4953f
C199 comp_p_5/vinn comp_p_5/latch_right 0.00802f
C200 vin comp_p_3/vinn 0.65736f
C201 vdd comp_p_6/latch_right 1.95583f
C202 comp_p_1/vinn vdd 1.45676f
C203 d2 comp_p_1/tail 0
C204 d4 comp_p_3/tail 0
C205 d4 d3 2.89503f
C206 d1 d3 0.32128f
C207 comp_p_6/vbias_p d3 0
C208 vin d2 0.72189f
C209 comp_p_5/vinn d6 0.00479f
C210 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vdd 0
C211 comp_p_2/latch_right comp_p_3/vinn 0.17373f
C212 d5 comp_p_3/out_left 0.02324f
C213 comp_p_1/vinn comp_p_0/vinn 0.94536f
C214 d5 vdd 2.4762f
C215 d4 comp_p_1/tail 0
C216 d1 comp_p_1/tail 0.00454f
C217 comp_p_6/vinn comp_p_4/latch_left 0.00606f
C218 comp_p_0/latch_left comp_p_2/out_left 0.01472f
C219 d4 vin 0.74069f
C220 vin d1 0.63586f
C221 comp_p_2/latch_right d2 0.00137f
C222 vin comp_p_6/vbias_p 1.44181f
C223 d4 comp_p_4/latch_right 0
C224 comp_p_6/vbias_p comp_p_4/latch_right 0.40389f
C225 d4 comp_p_6/tail 0.00252f
C226 comp_p_5/out_left comp_p_4/tail 0
C227 comp_p_2/latch_right d1 0.01472f
C228 comp_p_3/vinn comp_p_2/vinn 0.31181f
C229 comp_p_2/latch_right comp_p_6/vbias_p 0.39369f
C230 d3 comp_p_1/tail 0
C231 tmux_7therm_to_3bin_0/buffer_0/out d6 0
C232 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin tmux_7therm_to_3bin_0/R1/R1 0
C233 comp_p_3/tail vin 0.00233f
C234 vin d3 0.00158f
C235 d5 comp_p_1/vinn 0
C236 vbias_generation_0/XR_bias_2/R2 comp_p_6/vinn 0.00358f
C237 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vdd 0.00186f
C238 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin vdd 0.00196f
C239 d4 tmux_7therm_to_3bin_0/buffer_4/out 0
C240 comp_p_4/out_left vdd 0.02489f
C241 d5 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin 0.00355f
C242 comp_p_1/out_left comp_p_0/tail 0
C243 vin comp_p_1/tail 0.00233f
C244 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d4 0.00285f
C245 comp_p_6/vbias_p comp_p_2/vinn 0.12413f
C246 comp_p_1/latch_right d2 0.00123f
C247 comp_p_1/latch_left d6 0
C248 d4 comp_p_6/out_left 0.27385f
C249 tmux_7therm_to_3bin_0/R1/m1_n100_n100# d3 0
C250 comp_p_6/out_left comp_p_6/vbias_p -0.05282f
C251 vin comp_p_4/latch_right 0.21628f
C252 comp_p_5/vinn vdd 1.45079f
C253 d2 tmux_7therm_to_3bin_0/buffer_2/out 0
C254 vin comp_p_6/tail 0
C255 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin d6 0
C256 comp_p_2/latch_right vin 0.21614f
C257 comp_p_5/out_left d6 0
C258 d4 comp_p_1/latch_right 0.00137f
C259 comp_p_1/latch_right d1 0.09485f
C260 d0 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C261 comp_p_3/latch_left d6 0
C262 d1 tmux_7therm_to_3bin_0/buffer_2/out 0.00646f
C263 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d3 0
C264 comp_p_5/tail d6 0
C265 d2 tmux_7therm_to_3bin_0/R1/R1 0.00771f
C266 comp_p_0/latch_right d2 0.01472f
C267 d5 tmux_7therm_to_3bin_0/buffer_5/out 0
C268 comp_p_3/latch_right d6 0.00265f
C269 d5 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin 0
C270 d5 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin 0
C271 comp_p_4/latch_left vdd 0
C272 d4 tmux_7therm_to_3bin_0/R1/R1 0
C273 comp_p_1/latch_right d3 0
C274 d1 tmux_7therm_to_3bin_0/R1/R1 0.01255f
C275 comp_p_0/latch_right d1 0
C276 vin comp_p_2/vinn 0.52215f
C277 comp_p_0/latch_right comp_p_6/vbias_p 0.40389f
C278 tmux_7therm_to_3bin_0/buffer_0/out vdd 0
C279 dout0 dout1 -0
C280 comp_p_6/out_left vin 0.06197f
C281 comp_p_2/latch_right comp_p_2/vinn 0
C282 comp_p_0/latch_left comp_p_6/vbias_p 0.37827f
C283 comp_p_1/out_left d2 0
C284 d4 vbias_generation_0/bias_n 0.00802f
C285 comp_p_6/vbias_p vbias_generation_0/bias_n 0
C286 comp_p_1/latch_left vdd 2.04615f
C287 d3 tmux_7therm_to_3bin_0/R1/R1 0
C288 d2 d0 0.03267f
C289 comp_p_1/out_left d4 0
C290 comp_p_1/out_left d1 0.67001f
C291 comp_p_1/out_left comp_p_6/vbias_p -0.065f
C292 comp_p_3/out_left comp_p_5/out_left 0.01584f
C293 vdd comp_p_5/out_left 1.8042f
C294 d4 d0 0.03813f
C295 d1 d0 1.08821f
C296 comp_p_6/vbias_p d0 0.00463f
C297 comp_p_0/latch_right vin 0.21598f
C298 vdd tmux_7therm_to_3bin_0/buffer_7/in 0.0027f
C299 comp_p_2/latch_left comp_p_3/vinn 0.15294f
C300 comp_p_3/latch_left vdd 2.03617f
C301 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin d6 0
C302 vdd comp_p_5/tail 0.35567f
C303 d5 tmux_7therm_to_3bin_0/buffer_0/out 0
C304 comp_p_3/latch_right vdd 1.95376f
C305 comp_p_1/out_left d3 0
C306 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vdd 0
C307 comp_p_0/latch_left vin 0.00334f
C308 comp_p_0/latch_right comp_p_2/latch_right 0.01494f
C309 comp_p_5/vinn comp_p_4/out_left 0.01843f
C310 comp_p_0/out_left comp_p_2/out_left 0.09264f
C311 comp_p_1/vinn comp_p_1/latch_left 0.0067f
C312 vbias_generation_0/XR_bias_4/R1 comp_p_6/vbias_p 0.02724f
C313 vin vbias_generation_0/bias_n 0.0214f
C314 d3 d0 0.0327f
C315 d4 comp_p_4/tail -0.00224f
C316 comp_p_6/vbias_p comp_p_4/tail 0.31443f
C317 d4 comp_p_6/latch_left 0.06068f
C318 comp_p_4/vinn vdd 0.03662f
C319 comp_p_4/latch_right vbias_generation_0/bias_n 0
C320 comp_p_1/out_left vin 0.07139f
C321 d5 comp_p_1/latch_left 0
C322 comp_p_2/out_left vdd 0.02487f
C323 comp_p_2/latch_left comp_p_6/vbias_p 0.37827f
C324 d4 comp_p_5/latch_left 0.06548f
C325 comp_p_3/vinn d6 0
C326 d5 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin 0
C327 comp_p_2/tail comp_p_3/vinn 0.14685f
C328 comp_p_2/out_left comp_p_0/vinn 0.0271f
C329 d5 comp_p_5/out_left 0
C330 d4 comp_p_6/vinn 0.06841f
C331 comp_p_6/vbias_p comp_p_6/vinn 0.31983f
C332 tmux_7therm_to_3bin_0/buffer_6/out d6 0
C333 d4 comp_p_5/latch_right 0.06583f
C334 d5 comp_p_3/latch_left 0
C335 comp_p_0/tail vdd 0.00166f
C336 d2 d6 0.0531f
C337 comp_p_2/tail d2 -0.00224f
C338 d5 comp_p_3/latch_right 0.00185f
C339 vbias_generation_0/XR_bias_4/R1 vin 0.00472f
C340 comp_p_5/vinn comp_p_4/latch_left 0.16266f
C341 vin comp_p_4/tail 0.01181f
C342 d4 d6 0.76607f
C343 comp_p_1/vinn comp_p_2/out_left 0.00265f
C344 tmux_7therm_to_3bin_0/buffer_2/out tmux_7therm_to_3bin_0/R1/R1 0
C345 d1 d6 0.06436f
C346 comp_p_6/out_left vbias_generation_0/bias_n 0.00925f
C347 d4 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0
C348 vbias_generation_0/XR_bias_4/R1 comp_p_4/latch_right 0
C349 vin comp_p_6/latch_left 0.00266f
C350 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vdd 0
C351 comp_p_2/tail comp_p_6/vbias_p 0.31443f
C352 comp_p_2/latch_left vin 0.00664f
C353 comp_p_5/latch_left comp_p_4/latch_right 0.02598f
C354 vin comp_p_6/vinn 1.01745f
C355 comp_p_1/vinn comp_p_0/tail 0.10698f
C356 comp_p_3/tail d6 0
C357 d3 d6 0.07956f
C358 d3 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin 0.00238f
C359 comp_p_4/latch_right comp_p_6/vinn 0.00583f
C360 tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G d1 0
C361 comp_p_3/vinn comp_p_3/out_left 0.20126f
C362 comp_p_1/tail d6 0
C363 comp_p_5/vinn comp_p_5/out_left 0.19629f
C364 comp_p_3/vinn vdd 1.48772f
C365 vin d6 0.01178f
C366 comp_p_2/tail vin 0.0104f
C367 comp_p_1/out_left comp_p_0/latch_right 0
C368 comp_p_2/latch_left comp_p_2/vinn 0
C369 comp_p_3/vinn comp_p_0/vinn 0.53348f
C370 d2 comp_p_3/out_left 0.67197f
C371 comp_p_4/out_left comp_p_4/vinn 0.02516f
C372 d5 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin 0
C373 d2 vdd 1.1604f
C374 comp_p_0/out_left comp_p_6/vbias_p 0.68478f
C375 comp_p_2/out_left comp_p_4/out_left 0.01584f
C376 d0 tmux_7therm_to_3bin_0/R1/R1 0.00538f
C377 d4 comp_p_3/out_left 0.00143f
C378 d4 vdd 1.47711f
C379 d1 vdd 1.17278f
C380 comp_p_6/vbias_p comp_p_3/out_left -0.06014f
C381 comp_p_6/vbias_p vdd 12.48415f
C382 comp_p_5/vinn comp_p_4/vinn 0.32186f
C383 comp_p_6/out_left comp_p_6/vinn 0.14972f
C384 comp_p_1/vinn comp_p_3/vinn 0.03321f
C385 d1 comp_p_0/vinn -0
C386 tmux_7therm_to_3bin_0/buffer_4/out d6 0
C387 comp_p_6/vbias_p comp_p_0/vinn 0.12306f
C388 d5 comp_p_3/vinn 0
C389 comp_p_2/tail comp_p_2/vinn 0
C390 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin d6 0
C391 comp_p_1/vinn d2 0.00152f
C392 comp_p_1/out_left d0 -0
C393 comp_p_3/tail vdd 0.35691f
C394 d3 vdd 2.36726f
C395 d6.t1 vss 0.09613f
C396 d6.t0 vss 0.09121f
C397 d6.n0 vss 0.27214f
C398 d6.n1 vss 2.91721f
C399 d6.n2 vss 2.98722f
C400 comp_p_6/out_left.t1 vss 0.35725f
C401 comp_p_6/out_left.n0 vss 0.35824f
C402 comp_p_6/out_left.t2 vss 0.95164f
C403 comp_p_6/out_left.n1 vss 1.72525f
C404 comp_p_6/out_left.t0 vss 0.94389f
C405 comp_p_6/out_left.n2 vss 0.3128f
C406 comp_p_6/out_left.n3 vss 1.23781f
C407 d5.t0 vss 0.12676f
C408 d5.t1 vss 0.13359f
C409 d5.n0 vss 0.3782f
C410 d5.n1 vss 1.56109f
C411 d5.n2 vss 0.56227f
C412 d5.n3 vss 17.5754f
C413 comp_p_5/latch_right.t1 vss 0.4606f
C414 comp_p_5/latch_right.n0 vss 0.90852f
C415 comp_p_5/latch_right.t3 vss 1.93136f
C416 comp_p_5/latch_right.t2 vss 1.7936f
C417 comp_p_5/latch_right.n1 vss 3.06813f
C418 comp_p_5/latch_right.t0 vss 1.53795f
C419 comp_p_5/latch_right.n2 vss 0.44996f
C420 comp_p_5/latch_right.n3 vss 2.026f
C421 comp_p_5/latch_right.n4 vss 0.28331f
C422 comp_p_5/latch_left.t0 vss 1.25281f
C423 comp_p_5/latch_left.t3 vss 1.57061f
C424 comp_p_5/latch_left.t2 vss 1.45859f
C425 comp_p_5/latch_left.n0 vss 2.77309f
C426 comp_p_5/latch_left.n1 vss 1.77973f
C427 comp_p_5/latch_left.t1 vss 0.37457f
C428 comp_p_5/latch_left.n2 vss 1.60078f
C429 d4.t1 vss 0.07083f
C430 d4.t0 vss 0.06721f
C431 d4.n0 vss 0.20053f
C432 d4.n1 vss 4.3116f
C433 d4.n2 vss 6.94368f
C434 comp_p_4/out_left.t1 vss 0.26539f
C435 comp_p_4/out_left.n0 vss 0.26612f
C436 comp_p_4/out_left.t2 vss 0.70693f
C437 comp_p_4/out_left.n1 vss 1.28162f
C438 comp_p_4/out_left.t0 vss 0.70117f
C439 comp_p_4/out_left.n2 vss 0.23237f
C440 comp_p_4/out_left.n3 vss 0.91952f
C441 d3.t0 vss 0.10595f
C442 d3.t1 vss 0.11166f
C443 d3.n0 vss 0.31612f
C444 d3.n1 vss 2.45175f
C445 d3.n2 vss 0.37794f
C446 d3.n3 vss 6.98756f
C447 comp_p_3/latch_left.t0 vss 1.25281f
C448 comp_p_3/latch_left.t3 vss 1.57061f
C449 comp_p_3/latch_left.t2 vss 1.45859f
C450 comp_p_3/latch_left.n0 vss 2.77309f
C451 comp_p_3/latch_left.n1 vss 1.77973f
C452 comp_p_3/latch_left.t1 vss 0.37457f
C453 comp_p_3/latch_left.n2 vss 1.60078f
C454 d2.t1 vss 0.08704f
C455 d2.t0 vss 0.08259f
C456 d2.n0 vss 0.24464f
C457 d2.n1 vss 0.05352f
C458 d2.n2 vss 3.12412f
C459 d2.n3 vss 0.17713f
C460 d2.n4 vss 6.65299f
C461 comp_p_2/out_left.t1 vss 0.26539f
C462 comp_p_2/out_left.n0 vss 0.26612f
C463 comp_p_2/out_left.t2 vss 0.70693f
C464 comp_p_2/out_left.n1 vss 1.28162f
C465 comp_p_2/out_left.t0 vss 0.70117f
C466 comp_p_2/out_left.n2 vss 0.23237f
C467 comp_p_2/out_left.n3 vss 0.91952f
C468 comp_p_2/latch_left.t0 vss 1.01079f
C469 comp_p_2/latch_left.t3 vss 1.2672f
C470 comp_p_2/latch_left.t2 vss 1.17681f
C471 comp_p_2/latch_left.n0 vss 2.23738f
C472 comp_p_2/latch_left.n1 vss 1.43592f
C473 comp_p_2/latch_left.t1 vss 0.30221f
C474 comp_p_2/latch_left.n2 vss 1.29154f
C475 d1.t0 vss 0.06253f
C476 d1.t1 vss 0.0659f
C477 d1.n0 vss 0.18658f
C478 d1.n1 vss 2.95125f
C479 d1.n2 vss 1.63556f
C480 comp_p_0/out_left.t1 vss 0.26539f
C481 comp_p_0/out_left.n0 vss 0.26612f
C482 comp_p_0/out_left.t2 vss 0.70693f
C483 comp_p_0/out_left.n1 vss 1.28162f
C484 comp_p_0/out_left.t0 vss 0.70117f
C485 comp_p_0/out_left.n2 vss 0.23237f
C486 comp_p_0/out_left.n3 vss 0.91952f
C487 comp_p_0/latch_right.t1 vss 0.38673f
C488 comp_p_0/latch_right.n0 vss 0.76282f
C489 comp_p_0/latch_right.t3 vss 1.62161f
C490 comp_p_0/latch_right.t2 vss 1.50595f
C491 comp_p_0/latch_right.n1 vss 2.57607f
C492 comp_p_0/latch_right.t0 vss 1.2913f
C493 comp_p_0/latch_right.n2 vss 0.3778f
C494 comp_p_0/latch_right.n3 vss 1.70107f
C495 comp_p_0/latch_right.n4 vss 0.23787f
C496 vin.t4 vss 0.59408f
C497 vin.t5 vss 0.59368f
C498 vin.n0 vss 0.79767f
C499 vin.n1 vss 0.6245f
C500 vin.t6 vss 0.44152f
C501 vin.n2 vss 0.71826f
C502 vin.t7 vss 0.44095f
C503 vin.n3 vss 0.70618f
C504 vin.n4 vss 0.3347f
C505 vin.t8 vss 0.59408f
C506 vin.t9 vss 0.59368f
C507 vin.n5 vss 0.79767f
C508 vin.n6 vss 0.6245f
C509 vin.t10 vss 0.44152f
C510 vin.n7 vss 0.71826f
C511 vin.t11 vss 0.44095f
C512 vin.n8 vss 0.70618f
C513 vin.n9 vss 0.3347f
C514 vin.n10 vss 4.91504f
C515 vin.t16 vss 0.59408f
C516 vin.t17 vss 0.59368f
C517 vin.n11 vss 0.79767f
C518 vin.n12 vss 0.6245f
C519 vin.t18 vss 0.44152f
C520 vin.n13 vss 0.71826f
C521 vin.t19 vss 0.44095f
C522 vin.n14 vss 0.70618f
C523 vin.n15 vss 0.3347f
C524 vin.n16 vss 2.8404f
C525 vin.n17 vss 1.64812f
C526 vin.t24 vss 0.59408f
C527 vin.t25 vss 0.59368f
C528 vin.n18 vss 0.79767f
C529 vin.n19 vss 0.6245f
C530 vin.t26 vss 0.44152f
C531 vin.n20 vss 0.71826f
C532 vin.t27 vss 0.44095f
C533 vin.n21 vss 0.70618f
C534 vin.n22 vss 0.3347f
C535 vin.t0 vss 0.59408f
C536 vin.t1 vss 0.59368f
C537 vin.n23 vss 0.79767f
C538 vin.n24 vss 0.6245f
C539 vin.t2 vss 0.44152f
C540 vin.n25 vss 0.71826f
C541 vin.t3 vss 0.44095f
C542 vin.n26 vss 0.70618f
C543 vin.n27 vss 0.3239f
C544 vin.n28 vss 1.52012f
C545 vin.t12 vss 0.59408f
C546 vin.t13 vss 0.59368f
C547 vin.n29 vss 0.79767f
C548 vin.n30 vss 0.6245f
C549 vin.t14 vss 0.44152f
C550 vin.n31 vss 0.71826f
C551 vin.t15 vss 0.44095f
C552 vin.n32 vss 0.70618f
C553 vin.n33 vss 0.3329f
C554 vin.n34 vss 0.34148f
C555 vin.n35 vss 5.07332f
C556 vin.t20 vss 0.59408f
C557 vin.t21 vss 0.59368f
C558 vin.n36 vss 0.79767f
C559 vin.n37 vss 0.6245f
C560 vin.t22 vss 0.44152f
C561 vin.n38 vss 0.71826f
C562 vin.t23 vss 0.44095f
C563 vin.n39 vss 0.70618f
C564 vin.n40 vss 0.32699f
C565 vin.n41 vss 0.44314f
C566 vin.n42 vss 3.94534f
C567 vin.n43 vss 3.63034f
C568 vin.n44 vss 1.93785f
C569 vin.n45 vss 1.86451f
C570 d0.t1 vss 0.07748f
C571 d0.t0 vss 0.07351f
C572 d0.n0 vss 0.21724f
C573 d0.n1 vss 0.0497f
C574 d0.n2 vss 1.17415f
C575 d0.n3 vss 0.92124f
C576 comp_p_1/latch_left.t0 vss 1.25281f
C577 comp_p_1/latch_left.t3 vss 1.57061f
C578 comp_p_1/latch_left.t2 vss 1.45859f
C579 comp_p_1/latch_left.n0 vss 2.77309f
C580 comp_p_1/latch_left.n1 vss 1.77973f
C581 comp_p_1/latch_left.t1 vss 0.37457f
C582 comp_p_1/latch_left.n2 vss 1.60078f
C583 vdd.n0 vss 2.61721f
C584 vdd.n1 vss 0.35756f
C585 vdd.n2 vss 0.26019f
C586 vdd.n3 vss 0.35275f
C587 vdd.n4 vss 0.06624f
C588 vdd.n5 vss 0.41954f
C589 vdd.n6 vss 0.54535f
C590 vdd.n7 vss 0.02162f
C591 vdd.n8 vss 0.14181f
C592 vdd.n9 vss 0.0391f
C593 vdd.n10 vss 0.021f
C594 vdd.n11 vss 1.38167f
C595 vdd.n12 vss 0.0524f
C596 vdd.n13 vss 0.05055f
C597 vdd.n14 vss 0.96493f
C598 vdd.n15 vss 0.05036f
C599 vdd.n16 vss 1.21125f
C600 vdd.n17 vss 0.35311f
C601 vdd.n18 vss 0.13112f
C602 vdd.n19 vss 1.10198f
C603 vdd.n20 vss 0.75786f
C604 vdd.n21 vss 0.22854f
C605 vdd.n22 vss 0.79838f
C606 vdd.n23 vss 0.29909f
C607 vdd.n24 vss 0.04644f
C608 vdd.n25 vss 0.05036f
C609 vdd.n26 vss 0.06025f
C610 vdd.n27 vss 0.04646f
C611 vdd.n28 vss 1.10897f
C612 vdd.n29 vss 1.56207f
C613 vdd.n30 vss 0.44362f
C614 vdd.n31 vss 0.1174f
C615 vdd.n32 vss 0.16204f
C616 vdd.n33 vss 0.03922f
C617 vdd.n34 vss 0.03621f
C618 vdd.n35 vss 0.27064f
C619 vdd.n36 vss 0.81257f
C620 vdd.n37 vss 0.25756f
C621 vdd.n38 vss 1.57746f
C622 vdd.n39 vss 0.05055f
C623 vdd.n40 vss 0.05055f
C624 vdd.n41 vss 0.83194f
C625 vdd.n42 vss 0.04646f
C626 vdd.n43 vss 0.14146f
C627 vdd.n44 vss 0.05036f
C628 vdd.n45 vss 0.05036f
C629 vdd.n46 vss 1.35091f
C630 vdd.n47 vss 1.58445f
C631 vdd.n48 vss 0.0391f
C632 vdd.n49 vss 0.0391f
C633 vdd.n50 vss 0.02162f
C634 vdd.n51 vss -0.10021f
C635 vdd.n52 vss 0.05065f
C636 vdd.n53 vss 0.05148f
C637 vdd.n54 vss 0.02373f
C638 vdd.n55 vss 1.2119f
C639 vdd.n56 vss 1.10897f
C640 vdd.n57 vss 0.05053f
C641 vdd.n58 vss 0.13764f
C642 vdd.n59 vss 0.03922f
C643 vdd.n60 vss 1.64806f
C644 vdd.n61 vss 0.0442f
C645 vdd.n62 vss 0.27064f
C646 vdd.n63 vss 0.44362f
C647 vdd.n64 vss 0.81257f
C648 vdd.n65 vss 0.25756f
C649 vdd.n66 vss 0.03621f
C650 vdd.n67 vss 0.03922f
C651 vdd.n68 vss 1.56207f
C652 vdd.n69 vss 0.31046f
C653 vdd.n70 vss 0.05053f
C654 vdd.n71 vss 0.13204f
C655 vdd.n72 vss 0.13112f
C656 vdd.n73 vss 0.05065f
C657 vdd.n74 vss 0.24893f
C658 vdd.n75 vss 1.11737f
C659 vdd.n76 vss 0.05148f
C660 vdd.n77 vss 0.45766f
C661 vdd.n78 vss 0.00716f
C662 vdd.n79 vss 0.14273f
C663 vdd.n80 vss 0.03922f
C664 vdd.n81 vss 4.66263f
C665 vdd.n82 vss 0.14183f
C666 vdd.n83 vss 0.00288f
C667 vdd.n84 vss 0.01265f
C668 vdd.n85 vss 0.01876f
C669 vdd.n86 vss 0.01205f
C670 vdd.n87 vss 0.01876f
C671 vdd.n88 vss 0.14113f
C672 vdd.n89 vss 0.01265f
C673 vdd.n90 vss 0.01205f
C674 vdd.n91 vss 0.01205f
C675 vdd.n92 vss 0.01205f
C676 vdd.n93 vss 0.14113f
C677 vdd.n94 vss 0.01247f
C678 vdd.n95 vss 0.01247f
C679 vdd.n96 vss 0.14113f
C680 vdd.n97 vss 0.01922f
C681 vdd.n98 vss 0.01922f
C682 vdd.n99 vss 0.00671f
C683 vdd.n100 vss 0.00963f
C684 vdd.n101 vss 0.15461f
C685 vdd.n102 vss 0.01922f
C686 vdd.n103 vss 0.01922f
C687 vdd.n104 vss 0.08979f
C688 vdd.n105 vss 0.05335f
C689 vdd.n106 vss 0.17302f
C690 vdd.n107 vss 0.00945f
C691 vdd.n108 vss 0.00963f
C692 vdd.n110 vss 0.12318f
C693 vdd.n111 vss 0.01876f
C694 vdd.n112 vss 0.01874f
C695 vdd.n113 vss 0.01876f
C696 vdd.n114 vss 0.11701f
C697 vdd.n115 vss 0.11701f
C698 vdd.n116 vss 0.01876f
C699 vdd.n117 vss 0.01876f
C700 vdd.n118 vss 0.01874f
C701 vdd.n119 vss 0.01876f
C702 vdd.n120 vss 0.58863f
C703 vdd.n121 vss 0.14113f
C704 vdd.n122 vss 0.58863f
C705 vdd.n123 vss 0.01876f
C706 vdd.n124 vss 0.01876f
C707 vdd.n125 vss 0.01247f
C708 vdd.n126 vss 0.01205f
C709 vdd.n127 vss 0.01265f
C710 vdd.n128 vss 0.01265f
C711 vdd.n129 vss 0.01205f
C712 vdd.n130 vss 0.00573f
C713 vdd.n131 vss 0.14113f
C714 vdd.n132 vss 0.00573f
C715 vdd.n133 vss 0.01205f
C716 vdd.n134 vss 0.01247f
C717 vdd.n135 vss 0.14113f
C718 vdd.n136 vss 0.01922f
C719 vdd.n137 vss 0.01922f
C720 vdd.n138 vss 0.00963f
C721 vdd.n139 vss 0.00671f
C722 vdd.n140 vss 0.15461f
C723 vdd.n141 vss 0.01922f
C724 vdd.n142 vss 0.01922f
C725 vdd.n143 vss 0.00963f
C726 vdd.n144 vss 0.05365f
C727 vdd.n145 vss 0.08979f
C728 vdd.n146 vss 0.08979f
C729 vdd.n147 vss 0.05335f
C730 vdd.n148 vss 0.00671f
C731 vdd.n150 vss 0.12318f
C732 vdd.n151 vss 0.01874f
C733 vdd.n152 vss 0.01876f
C734 vdd.n153 vss 0.01876f
C735 vdd.n154 vss 0.11701f
C736 vdd.n155 vss 0.11701f
C737 vdd.n156 vss 0.01876f
C738 vdd.n157 vss 0.01874f
C739 vdd.n158 vss 0.01876f
C740 vdd.n159 vss 0.01876f
C741 vdd.n160 vss 0.1179f
C742 vdd.n161 vss 0.1179f
C743 vdd.n162 vss 0.14113f
C744 vdd.n163 vss 0.01247f
C745 vdd.n164 vss 0.01247f
C746 vdd.n165 vss 0.01203f
C747 vdd.n166 vss 0.00286f
C748 vdd.n167 vss 0.14968f
C749 vdd.n168 vss 0.55152f
C750 vdd.n169 vss 0.94598f
C751 vdd.n170 vss 0.00286f
C752 vdd.n171 vss 0.16815f
C753 vdd.n172 vss 0.00288f
C754 vdd.n173 vss 0.01265f
C755 vdd.n174 vss 0.01876f
C756 vdd.n175 vss 0.01205f
C757 vdd.n176 vss 0.01876f
C758 vdd.n177 vss 0.28226f
C759 vdd.n178 vss 0.01247f
C760 vdd.n179 vss 0.01876f
C761 vdd.n180 vss 0.28226f
C762 vdd.n181 vss 0.01922f
C763 vdd.n182 vss 0.01922f
C764 vdd.n183 vss 0.01874f
C765 vdd.n184 vss 0.00671f
C766 vdd.n185 vss 0.00671f
C767 vdd.n186 vss 0.13347f
C768 vdd.n187 vss 0.00963f
C769 vdd.n188 vss 0.01922f
C770 vdd.n189 vss 0.01922f
C771 vdd.n190 vss 0.28226f
C772 vdd.n191 vss 0.01922f
C773 vdd.n192 vss 0.01922f
C774 vdd.n193 vss 0.00963f
C775 vdd.n194 vss 0.01922f
C776 vdd.n195 vss 0.01922f
C777 vdd.n196 vss 0.00963f
C778 vdd.n197 vss 0.01876f
C779 vdd.n198 vss 0.01874f
C780 vdd.n199 vss 0.01876f
C781 vdd.n200 vss 0.01876f
C782 vdd.n201 vss 0.23402f
C783 vdd.n202 vss 0.01876f
C784 vdd.n203 vss 0.01876f
C785 vdd.n204 vss 0.23402f
C786 vdd.n205 vss 0.01876f
C787 vdd.n206 vss 0.01876f
C788 vdd.n207 vss 0.01874f
C789 vdd.n208 vss 0.01876f
C790 vdd.n209 vss 0.23581f
C791 vdd.n210 vss 0.01876f
C792 vdd.n211 vss 0.01874f
C793 vdd.n212 vss 0.00671f
C794 vdd.n213 vss 0.02985f
C795 vdd.n214 vss 0.13347f
C796 vdd.n215 vss 0.03002f
C797 vdd.n216 vss 0.00671f
C798 vdd.n217 vss 0.00963f
C799 vdd.n218 vss 0.01876f
C800 vdd.n219 vss 0.01876f
C801 vdd.n220 vss 0.23581f
C802 vdd.n221 vss 0.23581f
C803 vdd.n222 vss 0.01247f
C804 vdd.n223 vss 0.01265f
C805 vdd.n224 vss 0.01205f
C806 vdd.n225 vss 0.01205f
C807 vdd.n226 vss 0.01205f
C808 vdd.n227 vss 0.28226f
C809 vdd.n228 vss 0.00573f
C810 vdd.n229 vss 0.00573f
C811 vdd.n230 vss 0.01205f
C812 vdd.n231 vss 0.01205f
C813 vdd.n232 vss 0.01247f
C814 vdd.n233 vss 0.01205f
C815 vdd.n234 vss 0.01265f
C816 vdd.n235 vss 0.01265f
C817 vdd.n236 vss 0.01203f
C818 vdd.n237 vss 0.01247f
C819 vdd.n238 vss 0.01876f
C820 vdd.n239 vss 0.01876f
C821 vdd.n240 vss 0.01205f
C822 vdd.n241 vss 0.01205f
C823 vdd.n242 vss 0.01876f
C824 vdd.n243 vss 0.01876f
C825 vdd.n244 vss 0.28226f
C826 vdd.n245 vss 0.01247f
C827 vdd.n246 vss 0.01247f
C828 vdd.n247 vss 0.01265f
C829 vdd.n248 vss 0.00288f
C830 vdd.n249 vss 0.00671f
C831 vdd.n250 vss 0.00963f
C832 vdd.n251 vss 0.01922f
C833 vdd.n252 vss 0.01922f
C834 vdd.n253 vss 0.28226f
C835 vdd.n254 vss 0.01922f
C836 vdd.n255 vss 0.01922f
C837 vdd.n256 vss 0.00963f
C838 vdd.n257 vss 0.28226f
C839 vdd.n258 vss 0.01876f
C840 vdd.n259 vss 0.01922f
C841 vdd.n260 vss 0.01922f
C842 vdd.n261 vss 0.00671f
C843 vdd.n262 vss 0.00963f
C844 vdd.n263 vss 0.01922f
C845 vdd.n264 vss 0.01922f
C846 vdd.n265 vss 0.01874f
C847 vdd.n266 vss 0.13347f
C848 vdd.n267 vss 0.04809f
C849 vdd.n268 vss 0.00671f
C850 vdd.n269 vss 0.00963f
C851 vdd.n270 vss 0.01876f
C852 vdd.n271 vss 0.01876f
C853 vdd.n272 vss 0.23581f
C854 vdd.n273 vss 0.01876f
C855 vdd.n274 vss 0.01876f
C856 vdd.n275 vss 0.01874f
C857 vdd.n276 vss 0.01876f
C858 vdd.n277 vss 0.23402f
C859 vdd.n278 vss 0.01876f
C860 vdd.n279 vss 0.01876f
C861 vdd.n280 vss 0.23402f
C862 vdd.n281 vss 0.01876f
C863 vdd.n282 vss 0.01876f
C864 vdd.n283 vss 0.01874f
C865 vdd.n284 vss 0.01876f
C866 vdd.n285 vss 0.28226f
C867 vdd.n286 vss 0.01247f
C868 vdd.n287 vss 0.01247f
C869 vdd.n288 vss 0.01205f
C870 vdd.n289 vss 0.01205f
C871 vdd.n290 vss 0.01205f
C872 vdd.n291 vss 0.00573f
C873 vdd.n292 vss 0.28226f
C874 vdd.n293 vss 0.01205f
C875 vdd.n294 vss 0.01265f
C876 vdd.n295 vss 0.01205f
C877 vdd.n296 vss 0.01205f
C878 vdd.n297 vss 0.00573f
C879 vdd.n298 vss 0.28226f
C880 vdd.n299 vss 0.28226f
C881 vdd.n300 vss 0.01265f
C882 vdd.n301 vss 0.01265f
C883 vdd.n302 vss 0.01205f
C884 vdd.n303 vss 0.01247f
C885 vdd.n304 vss 0.01876f
C886 vdd.n305 vss 0.01876f
C887 vdd.n306 vss 0.23581f
C888 vdd.n307 vss 0.23581f
C889 vdd.n308 vss 0.01876f
C890 vdd.n309 vss 0.01874f
C891 vdd.n310 vss 0.00671f
C892 vdd.n311 vss 0.02985f
C893 vdd.n312 vss 0.13347f
C894 vdd.n313 vss 0.1065f
C895 vdd.n314 vss 0.08433f
C896 vdd.n315 vss 0.00286f
C897 vdd.n316 vss 0.01203f
C898 vdd.n317 vss 0.01247f
C899 vdd.n318 vss 0.01876f
C900 vdd.n319 vss 0.01876f
C901 vdd.n320 vss 0.23581f
C902 vdd.n321 vss 0.23581f
C903 vdd.n322 vss 0.01247f
C904 vdd.n323 vss 0.01247f
C905 vdd.n324 vss 0.01876f
C906 vdd.n325 vss 0.01205f
C907 vdd.n326 vss 0.01265f
C908 vdd.n327 vss 0.01265f
C909 vdd.n328 vss 0.01205f
C910 vdd.n329 vss 0.01247f
C911 vdd.n330 vss 0.01876f
C912 vdd.n331 vss 0.01247f
C913 vdd.n332 vss 0.28226f
C914 vdd.n333 vss 0.01247f
C915 vdd.n334 vss 0.01205f
C916 vdd.n335 vss 0.01265f
C917 vdd.n336 vss 0.01265f
C918 vdd.n337 vss 0.01205f
C919 vdd.n338 vss 0.00288f
C920 vdd.n339 vss 0.00573f
C921 vdd.n340 vss 0.28226f
C922 vdd.n341 vss 0.00573f
C923 vdd.n342 vss 0.01205f
C924 vdd.n343 vss 0.01247f
C925 vdd.n344 vss 0.28226f
C926 vdd.n345 vss 0.01247f
C927 vdd.n346 vss 0.01247f
C928 vdd.n347 vss 0.01203f
C929 vdd.n348 vss 0.00286f
C930 vdd.n349 vss 0.08408f
C931 vdd.n350 vss 0.04502f
C932 vdd.n351 vss 0.61277f
C933 vdd.n352 vss 2.8122f
C934 vdd.n353 vss 0.00671f
C935 vdd.n354 vss 0.13347f
C936 vdd.n355 vss 0.00963f
C937 vdd.n356 vss 0.01922f
C938 vdd.n357 vss 0.01922f
C939 vdd.n358 vss 0.95388f
C940 vdd.n359 vss 0.01876f
C941 vdd.n360 vss 0.95388f
C942 vdd.n361 vss 0.01876f
C943 vdd.n362 vss 0.01876f
C944 vdd.n363 vss 0.01922f
C945 vdd.n364 vss 0.01922f
C946 vdd.n365 vss 0.01874f
C947 vdd.n366 vss 0.00963f
C948 vdd.n367 vss 0.01922f
C949 vdd.n368 vss 0.01922f
C950 vdd.n369 vss 0.95388f
C951 vdd.n370 vss 0.01876f
C952 vdd.n371 vss 0.01876f
C953 vdd.n372 vss 0.01876f
C954 vdd.n373 vss 0.95388f
C955 vdd.n374 vss 0.01922f
C956 vdd.n375 vss 0.01922f
C957 vdd.n376 vss 0.00963f
C958 vdd.n377 vss 0.01876f
C959 vdd.n378 vss 0.01874f
C960 vdd.n379 vss 0.01876f
C961 vdd.n380 vss 1.47933f
C962 vdd.n381 vss 0.01876f
C963 vdd.n382 vss 0.01874f
C964 vdd.n383 vss 0.00671f
C965 vdd.n384 vss 0.13347f
C966 vdd.n385 vss 0.02985f
C967 vdd.n386 vss 0.00671f
C968 vdd.n387 vss 0.00963f
C969 vdd.n388 vss 0.01876f
C970 vdd.n389 vss 0.01876f
C971 vdd.n390 vss 1.47933f
C972 vdd.n391 vss 0.01876f
C973 vdd.n392 vss 0.01874f
C974 vdd.n393 vss 0.00671f
C975 vdd.n394 vss 0.14448f
C976 vdd.n395 vss 0.7389f
C977 vdd.n396 vss 1.74058f
C978 vdd.n397 vss 0.00671f
C979 vdd.n398 vss 0.13347f
C980 vdd.n399 vss 0.00963f
C981 vdd.n400 vss 0.01922f
C982 vdd.n401 vss 0.01922f
C983 vdd.n402 vss 0.95388f
C984 vdd.n403 vss 0.01876f
C985 vdd.n404 vss 0.95388f
C986 vdd.n405 vss 0.01876f
C987 vdd.n406 vss 0.01876f
C988 vdd.n407 vss 0.01922f
C989 vdd.n408 vss 0.01922f
C990 vdd.n409 vss 0.01874f
C991 vdd.n410 vss 0.00963f
C992 vdd.n411 vss 0.01922f
C993 vdd.n412 vss 0.01922f
C994 vdd.n413 vss 0.95388f
C995 vdd.n414 vss 0.01876f
C996 vdd.n415 vss 0.01876f
C997 vdd.n416 vss 0.01876f
C998 vdd.n417 vss 0.95388f
C999 vdd.n418 vss 0.01922f
C1000 vdd.n419 vss 0.01922f
C1001 vdd.n420 vss 0.00963f
C1002 vdd.n421 vss 0.01876f
C1003 vdd.n422 vss 0.01874f
C1004 vdd.n423 vss 0.01876f
C1005 vdd.n424 vss 1.47933f
C1006 vdd.n425 vss 0.01876f
C1007 vdd.n426 vss 0.01874f
C1008 vdd.n427 vss 0.00671f
C1009 vdd.n428 vss 0.13347f
C1010 vdd.n429 vss 0.02985f
C1011 vdd.n430 vss 0.00671f
C1012 vdd.n431 vss 0.00963f
C1013 vdd.n432 vss 0.01876f
C1014 vdd.n433 vss 0.01876f
C1015 vdd.n434 vss 1.47933f
C1016 vdd.n435 vss 0.01876f
C1017 vdd.n436 vss 0.01874f
C1018 vdd.n437 vss 0.00671f
C1019 vdd.n438 vss 0.15087f
C1020 vdd.n439 vss 0.82136f
C1021 vdd.n440 vss 3.2949f
C1022 vdd.n441 vss 5.20887f
C1023 vdd.n442 vss 2.54816f
C1024 vdd.n443 vss 0.54302f
C1025 vdd.n444 vss 0.0175f
C1026 vdd.n445 vss 0.44678f
C1027 vdd.n446 vss 0.48198f
C1028 vdd.n447 vss 0.02162f
C1029 vdd.n448 vss 0.25976f
C1030 vdd.n449 vss 0.0391f
C1031 vdd.n450 vss 0.0442f
C1032 vdd.n451 vss 2.76335f
C1033 vdd.n452 vss 0.03922f
C1034 vdd.n453 vss 0.03922f
C1035 vdd.n454 vss 0.49785f
C1036 vdd.n455 vss 0.0391f
C1037 vdd.n456 vss 0.0442f
C1038 vdd.n457 vss 0.14273f
C1039 vdd.n458 vss -0.10021f
C1040 vdd.n459 vss 0.02162f
C1041 vdd.n460 vss 0.0442f
C1042 vdd.n461 vss 0.03621f
C1043 vdd.n462 vss 0.62091f
C1044 vdd.n463 vss 0.03922f
C1045 vdd.n464 vss 2.70181f
C1046 vdd.n465 vss 0.03922f
C1047 vdd.n466 vss 0.13204f
C1048 vdd.n467 vss 0.25756f
C1049 vdd.n468 vss 0.81257f
C1050 vdd.n469 vss 0.05065f
C1051 vdd.n470 vss 0.05065f
C1052 vdd.n471 vss 3.02905f
C1053 vdd.n472 vss 0.05065f
C1054 vdd.n473 vss 0.05065f
C1055 vdd.n474 vss 0.03621f
C1056 vdd.n475 vss 0.0442f
C1057 vdd.n476 vss 0.25756f
C1058 vdd.n477 vss 0.81257f
C1059 vdd.n478 vss 0.13204f
C1060 vdd.n479 vss 0.13112f
C1061 vdd.n480 vss 0.14146f
C1062 vdd.n481 vss 0.45766f
C1063 vdd.n482 vss 0.05036f
C1064 vdd.n483 vss 0.05055f
C1065 vdd.n484 vss 0.83194f
C1066 vdd.n485 vss 0.27215f
C1067 vdd.n486 vss 3.15491f
C1068 vdd.n487 vss 0.06025f
C1069 vdd.n488 vss 3.02905f
C1070 vdd.n489 vss 0.05053f
C1071 vdd.n490 vss 0.05053f
C1072 vdd.n491 vss 0.81257f
C1073 vdd.n492 vss 0.01837f
C1074 vdd.n493 vss 0.27215f
C1075 vdd.n494 vss 0.05036f
C1076 vdd.n495 vss 0.0605f
C1077 vdd.n496 vss 3.1689f
C1078 vdd.n497 vss 0.05055f
C1079 vdd.n498 vss 0.05055f
C1080 vdd.n499 vss 2.23473f
C1081 vdd.n500 vss 0.05036f
C1082 vdd.n501 vss 0.0605f
C1083 vdd.n502 vss 0.05036f
C1084 vdd.n503 vss 0.25976f
C1085 vdd.n504 vss 0.00716f
C1086 vdd.n505 vss 0.05065f
C1087 vdd.n506 vss 0.05148f
C1088 vdd.n507 vss -0.10021f
C1089 vdd.n508 vss 3.12415f
C1090 vdd.n509 vss 0.05065f
C1091 vdd.n510 vss 0.05036f
C1092 vdd.n511 vss 0.01837f
C1093 vdd.n512 vss 2.76335f
C1094 vdd.n513 vss 0.05148f
C1095 vdd.n514 vss 0.05148f
C1096 vdd.n515 vss 0.13764f
C1097 vdd.n516 vss 0.13139f
C1098 vdd.n517 vss 0.02162f
C1099 vdd.n518 vss 0.0391f
C1100 vdd.n519 vss 0.03922f
C1101 vdd.n520 vss 0.03621f
C1102 vdd.n521 vss 0.25756f
C1103 vdd.n522 vss 0.0442f
C1104 vdd.n523 vss 0.03922f
C1105 vdd.n524 vss 0.03922f
C1106 vdd.n525 vss 0.44362f
C1107 vdd.n526 vss 0.02373f
C1108 vdd.n527 vss 0.13204f
C1109 vdd.n528 vss 0.13112f
C1110 vdd.n529 vss 0.14146f
C1111 vdd.n530 vss 0.14273f
C1112 vdd.n531 vss 0.00716f
C1113 vdd.n532 vss 0.45766f
C1114 vdd.n533 vss 0.83194f
C1115 vdd.n534 vss 0.25976f
C1116 vdd.n535 vss 2.56756f
C1117 vdd.n536 vss 0.03922f
C1118 vdd.n537 vss 0.0391f
C1119 vdd.n538 vss 0.03621f
C1120 vdd.n539 vss 0.12836f
C1121 vdd.n540 vss 0.03922f
C1122 vdd.n541 vss 0.0442f
C1123 vdd.n542 vss 0.13204f
C1124 vdd.n543 vss 2.21795f
C1125 vdd.n544 vss 0.13112f
C1126 vdd.n545 vss 0.13139f
C1127 vdd.n546 vss 0.14273f
C1128 vdd.n547 vss 0.14146f
C1129 vdd.n548 vss 0.01837f
C1130 vdd.n549 vss 0.01837f
C1131 vdd.n550 vss 0.05036f
C1132 vdd.n551 vss 0.05053f
C1133 vdd.n552 vss 0.62091f
C1134 vdd.n553 vss 0.05053f
C1135 vdd.n554 vss 0.04646f
C1136 vdd.n555 vss 0.27064f
C1137 vdd.n556 vss 0.25756f
C1138 vdd.n557 vss 0.81257f
C1139 vdd.n558 vss 0.44362f
C1140 vdd.n559 vss 0.02373f
C1141 vdd.n560 vss 0.13764f
C1142 vdd.n561 vss 0.03922f
C1143 vdd.n562 vss 0.0391f
C1144 vdd.n563 vss 0.00819f
C1145 vdd.n564 vss 0.00819f
C1146 vdd.n565 vss 0.02162f
C1147 vdd.n566 vss 0.83967f
C1148 vdd.n567 vss 0.03616f
C1149 vdd.n568 vss 0.0175f
C1150 vdd.n569 vss 0.63687f
C1151 vdd.n570 vss 0.21822f
C1152 vdd.n571 vss 1.99771f
C1153 vdd.n572 vss 0.72869f
C1154 vdd.n573 vss 0.72409f
C1155 vdd.n574 vss 0.02162f
C1156 vdd.n575 vss 0.25976f
C1157 vdd.n576 vss 0.0391f
C1158 vdd.n577 vss 0.0442f
C1159 vdd.n578 vss 1.38167f
C1160 vdd.n579 vss 0.03922f
C1161 vdd.n580 vss 0.05055f
C1162 vdd.n581 vss 1.11737f
C1163 vdd.n582 vss 0.05036f
C1164 vdd.n583 vss 1.57746f
C1165 vdd.n584 vss 0.91019f
C1166 vdd.n585 vss 0.05065f
C1167 vdd.n586 vss 0.05065f
C1168 vdd.n587 vss 0.05066f
C1169 vdd.n589 vss 0.58501f
C1170 vdd.n590 vss 0.02897f
C1171 vdd.n591 vss 0.80577f
C1172 vdd.n592 vss 0.36203f
C1173 vdd.n593 vss 0.23995f
C1174 vdd.n594 vss 0.23661f
C1175 vdd.n595 vss 0.02867f
C1176 vdd.n596 vss 0.05287f
C1177 vdd.n597 vss 0.05148f
C1178 vdd.n598 vss 1.43602f
C1179 vdd.n599 vss 2.16166f
C1180 vdd.n600 vss 0.0605f
C1181 vdd.n601 vss 0.14273f
C1182 vdd.n602 vss 0.83194f
C1183 vdd.n603 vss 0.05065f
C1184 vdd.n604 vss 0.05148f
C1185 vdd.n605 vss -0.10021f
C1186 vdd.n606 vss 0.31046f
C1187 vdd.n607 vss 0.13139f
C1188 vdd.n608 vss 0.12836f
C1189 vdd.n609 vss 0.00819f
C1190 vdd.n610 vss 0.00819f
C1191 vdd.n611 vss 0.0391f
C1192 vdd.n612 vss 0.03922f
C1193 vdd.n613 vss 0.0442f
C1194 vdd.n614 vss 0.27064f
C1195 vdd.n615 vss 0.13112f
C1196 vdd.n616 vss 0.05036f
C1197 vdd.n617 vss 0.14146f
C1198 vdd.n618 vss 0.01837f
C1199 vdd.n619 vss 0.01837f
C1200 vdd.n620 vss 0.27215f
C1201 vdd.n621 vss 0.04644f
C1202 vdd.n622 vss 0.05036f
C1203 vdd.n623 vss 0.04646f
C1204 vdd.n624 vss 0.05053f
C1205 vdd.n625 vss 1.10897f
C1206 vdd.n626 vss 1.64806f
C1207 vdd.n627 vss 1.2119f
C1208 vdd.n628 vss 0.05053f
C1209 vdd.n629 vss 0.13204f
C1210 vdd.n630 vss 0.13764f
C1211 vdd.n631 vss 0.02373f
C1212 vdd.n632 vss 0.44362f
C1213 vdd.n633 vss 0.81257f
C1214 vdd.n634 vss 0.25756f
C1215 vdd.n635 vss 0.03621f
C1216 vdd.n636 vss 0.03922f
C1217 vdd.n637 vss 1.56207f
C1218 vdd.n638 vss 1.35091f
C1219 vdd.n639 vss 0.05065f
C1220 vdd.n640 vss 0.05148f
C1221 vdd.n641 vss 0.45766f
C1222 vdd.n642 vss 0.00716f
C1223 vdd.n643 vss 0.05055f
C1224 vdd.n644 vss 0.24893f
C1225 vdd.n645 vss 1.58445f
C1226 vdd.n646 vss 0.03922f
C1227 vdd.n647 vss 0.03616f
C1228 vdd.n648 vss 0.0175f
C1229 vdd.n649 vss 0.0387f
C1230 vdd.n650 vss 0.52082f
C1231 vdd.n651 vss 0.39448f
C1232 vdd.n652 vss 0.33684f
C1233 vdd.n653 vss 1.25827f
C1234 vdd.n654 vss 4.50133f
C1235 vdd.n655 vss 2.69174f
C1236 vdd.n656 vss 0.22837f
C1237 vdd.n657 vss 3.72504f
C1238 vdd.n658 vss 0.09923f
C1239 vdd.n659 vss 0.44678f
C1240 vdd.n660 vss 0.48198f
C1241 vdd.n661 vss 0.02884f
C1242 vdd.n662 vss 0.0175f
C1243 vdd.n663 vss 0.03616f
C1244 vdd.n664 vss 0.03922f
C1245 vdd.n665 vss 0.0442f
C1246 vdd.n666 vss 3.15491f
C1247 vdd.n667 vss 0.0442f
C1248 vdd.n668 vss 0.03922f
C1249 vdd.n669 vss 0.0391f
C1250 vdd.n670 vss 0.00819f
C1251 vdd.n671 vss 0.00819f
C1252 vdd.n672 vss 0.12836f
C1253 vdd.n673 vss -0.10021f
C1254 vdd.n674 vss 0.05065f
C1255 vdd.n675 vss 2.70181f
C1256 vdd.n676 vss 0.05065f
C1257 vdd.n677 vss 0.05148f
C1258 vdd.n678 vss 0.45766f
C1259 vdd.n679 vss 0.83194f
C1260 vdd.n680 vss 0.27215f
C1261 vdd.n681 vss 0.04644f
C1262 vdd.n682 vss 0.05055f
C1263 vdd.n683 vss 0.49785f
C1264 vdd.n684 vss 0.05055f
C1265 vdd.n685 vss 0.04644f
C1266 vdd.n686 vss 0.05036f
C1267 vdd.n687 vss 0.04646f
C1268 vdd.n688 vss 0.27064f
C1269 vdd.n689 vss 0.06025f
C1270 vdd.n690 vss 3.30035f
C1271 vdd.n691 vss 0.05055f
C1272 vdd.n692 vss 0.05055f
C1273 vdd.n693 vss 0.13112f
C1274 vdd.n694 vss 0.14146f
C1275 vdd.n695 vss 0.01837f
C1276 vdd.n696 vss 0.27064f
C1277 vdd.n697 vss 0.05053f
C1278 vdd.n698 vss 0.05053f
C1279 vdd.n699 vss 0.04644f
C1280 vdd.n700 vss 0.05036f
C1281 vdd.n701 vss 0.01837f
C1282 vdd.n702 vss 0.01837f
C1283 vdd.n703 vss 0.05036f
C1284 vdd.n704 vss 0.04646f
C1285 vdd.n705 vss 0.27064f
C1286 vdd.n706 vss 0.06025f
C1287 vdd.n707 vss 2.57036f
C1288 vdd.n708 vss 0.06025f
C1289 vdd.n709 vss 0.05053f
C1290 vdd.n710 vss 0.05036f
C1291 vdd.n711 vss 0.01837f
C1292 vdd.n712 vss 0.05036f
C1293 vdd.n713 vss 0.05053f
C1294 vdd.n714 vss 0.04646f
C1295 vdd.n715 vss 0.05036f
C1296 vdd.n716 vss 0.04644f
C1297 vdd.n717 vss 0.03616f
C1298 vdd.n718 vss 0.25976f
C1299 vdd.n719 vss 0.00716f
C1300 vdd.n720 vss 0.05148f
C1301 vdd.n721 vss 2.23473f
C1302 vdd.n722 vss 0.05148f
C1303 vdd.n723 vss 0.45766f
C1304 vdd.n724 vss 0.83194f
C1305 vdd.n725 vss 0.27215f
C1306 vdd.n726 vss 0.0605f
C1307 vdd.n727 vss 3.30315f
C1308 vdd.n728 vss 0.0605f
C1309 vdd.n729 vss 0.05055f
C1310 vdd.n730 vss 0.00716f
C1311 vdd.n731 vss 0.14273f
C1312 vdd.n732 vss 0.13139f
C1313 vdd.n733 vss 0.0391f
C1314 vdd.n734 vss 0.00819f
C1315 vdd.n735 vss 0.00819f
C1316 vdd.n736 vss 0.12836f
C1317 vdd.n737 vss -0.10021f
C1318 vdd.n738 vss 0.13764f
C1319 vdd.n739 vss 0.02373f
C1320 vdd.n740 vss 0.44362f
C1321 vdd.n741 vss 0.05148f
C1322 vdd.n742 vss 2.21795f
C1323 vdd.n743 vss 0.05148f
C1324 vdd.n744 vss 0.44362f
C1325 vdd.n745 vss 0.02373f
C1326 vdd.n746 vss 0.13764f
C1327 vdd.n747 vss 0.03922f
C1328 vdd.n748 vss 3.12415f
C1329 vdd.n749 vss 0.03922f
C1330 vdd.n750 vss 0.0391f
C1331 vdd.n751 vss 0.00819f
C1332 vdd.n752 vss 0.00819f
C1333 vdd.n753 vss 0.12836f
C1334 vdd.n754 vss 0.13139f
C1335 vdd.n755 vss 0.03922f
C1336 vdd.n756 vss 3.1689f
C1337 vdd.n757 vss 0.03922f
C1338 vdd.n758 vss 0.03616f
C1339 vdd.n759 vss 0.0175f
C1340 vdd.n760 vss 0.02884f
C1341 vdd.n761 vss 0.83967f
C1342 vdd.n762 vss 0.63703f
C1343 vdd.n763 vss 4.0112f
C1344 vdd.n764 vss 13.4668f
C1345 vdd.n765 vss 2.61946f
C1346 vdd.n766 vss 2.17473f
C1347 vdd.n767 vss 0.97899f
C1348 vdd.n768 vss 0.90949f
C1349 vdd.n769 vss 0.49844f
C1350 vdd.n770 vss 0.69134f
C1351 vdd.n771 vss 0.0535f
C1352 vdd.n772 vss 0.0175f
C1353 vdd.n773 vss 0.03616f
C1354 vdd.n774 vss 0.25976f
C1355 vdd.n775 vss 0.0442f
C1356 vdd.n776 vss 0.03922f
C1357 vdd.n777 vss 0.13139f
C1358 vdd.n778 vss 0.12836f
C1359 vdd.n779 vss 0.00819f
C1360 vdd.n780 vss 0.00819f
C1361 vdd.n781 vss 1.38167f
C1362 vdd.n782 vss 0.01837f
C1363 vdd.n783 vss 0.01837f
C1364 vdd.n784 vss 0.05036f
C1365 vdd.n785 vss 0.04644f
C1366 vdd.n786 vss 0.27215f
C1367 vdd.n787 vss 0.0605f
C1368 vdd.n788 vss 1.65158f
C1369 vdd.n789 vss 1.65018f
C1370 vdd.n790 vss 1.51453f
C1371 vdd.n791 vss 0.0442f
C1372 vdd.n792 vss 0.05148f
C1373 vdd.n793 vss 0.03486f
C1374 vdd.n794 vss 0.05031f
C1375 vdd.n795 vss 1.35091f
C1376 vdd.n796 vss 0.06718f
C1377 vdd.n797 vss 0.05958f
C1378 vdd.n798 vss 0.1284f
C1379 vdd.n799 vss 0.13085f
C1380 vdd.n800 vss 0.00819f
C1381 vdd.n801 vss 0.00819f
C1382 vdd.n802 vss 0.0391f
C1383 vdd.n803 vss 0.03922f
C1384 vdd.n804 vss 0.13413f
C1385 vdd.n805 vss 0.02373f
C1386 vdd.n806 vss 0.13204f
C1387 vdd.n807 vss 0.05053f
C1388 vdd.n808 vss 0.31046f
C1389 vdd.n809 vss 0.05053f
C1390 vdd.n810 vss 0.05036f
C1391 vdd.n811 vss 0.01837f
C1392 vdd.n812 vss 0.01837f
C1393 vdd.n813 vss 0.14146f
C1394 vdd.n814 vss 0.13492f
C1395 vdd.n815 vss 0.05248f
C1396 vdd.n816 vss 0.24893f
C1397 vdd.n817 vss 1.58445f
C1398 vdd.n818 vss 0.03673f
C1399 vdd.n819 vss 0.0358f
C1400 vdd.n820 vss 0.0175f
C1401 vdd.n821 vss 0.0535f
C1402 vdd.n822 vss 0.90949f
C1403 vdd.n823 vss 0.97899f
C1404 vdd.n824 vss 2.47098f
C1405 vdd.n825 vss 0.19252f
C1406 vdd.n826 vss 0.15002f
C1407 vdd.n827 vss 0.17331f
C1408 comp_p_6/vbias_p.t3 vss 0.68599f
C1409 comp_p_6/vbias_p.t2 vss 0.72093f
C1410 comp_p_6/vbias_p.n0 vss 1.08727f
C1411 comp_p_6/vbias_p.n1 vss 1.83582f
C1412 comp_p_6/vbias_p.t4 vss 0.68599f
C1413 comp_p_6/vbias_p.t6 vss 0.68599f
C1414 comp_p_6/vbias_p.t5 vss 0.68599f
C1415 comp_p_6/vbias_p.t7 vss 0.68599f
C1416 comp_p_6/vbias_p.n2 vss 2.59363f
C1417 comp_p_6/vbias_p.n3 vss 3.00042f
C1418 comp_p_6/vbias_p.n4 vss 0.8862f
C1419 comp_p_6/vbias_p.n5 vss 9.09667f
C1420 comp_p_6/vbias_p.n6 vss 0.28436f
C1421 comp_p_6/vbias_p.t0 vss 0.66669f
C1422 comp_p_6/vbias_p.t8 vss 0.72093f
C1423 comp_p_6/vbias_p.n7 vss 0.24364f
C1424 comp_p_6/vbias_p.n8 vss 1.2049f
C1425 comp_p_6/vbias_p.t1 vss 0.26392f
C1426 tmux_7therm_to_3bin_0/tmux_2to1_3/A vss 0.4939f
C1427 tmux_7therm_to_3bin_0/tmux_2to1_0/XM5/G vss 0.55051f
C1428 tmux_7therm_to_3bin_0/buffer_9/inv_1/vin vss 0.52606f
C1429 dout2 vss 0.32356f
C1430 tmux_7therm_to_3bin_0/buffer_8/inv_1/vin vss 0.52606f
C1431 dout1 vss 0.32356f
C1432 tmux_7therm_to_3bin_0/buffer_7/inv_1/vin vss 0.52606f
C1433 dout0 vss 0.32356f
C1434 tmux_7therm_to_3bin_0/buffer_6/inv_1/vin vss 0.5271f
C1435 tmux_7therm_to_3bin_0/buffer_6/out vss 0.64621f
C1436 d6 vss 10.21596f
C1437 tmux_7therm_to_3bin_0/buffer_5/inv_1/vin vss 0.52606f
C1438 tmux_7therm_to_3bin_0/buffer_5/out vss 0.6696f
C1439 d5 vss -3.15969f
C1440 vdd vss 0.37079p
C1441 tmux_7therm_to_3bin_0/buffer_4/inv_1/vin vss 0.52606f
C1442 tmux_7therm_to_3bin_0/buffer_4/out vss 0.70068f
C1443 d4 vss 8.90089f
C1444 tmux_7therm_to_3bin_0/buffer_3/inv_1/vin vss 0.52606f
C1445 tmux_7therm_to_3bin_0/R1/R2 vss 0.22083f
C1446 d3 vss 3.13204f
C1447 tmux_7therm_to_3bin_0/buffer_2/inv_1/vin vss 0.52811f
C1448 tmux_7therm_to_3bin_0/buffer_2/out vss 0.28552f
C1449 d2 vss 7.10238f
C1450 tmux_7therm_to_3bin_0/buffer_1/inv_1/vin vss 0.52606f
C1451 tmux_7therm_to_3bin_0/buffer_1/out vss 0.30295f
C1452 d1 vss 10.48549f
C1453 tmux_7therm_to_3bin_0/buffer_0/inv_1/vin vss 0.52606f
C1454 tmux_7therm_to_3bin_0/buffer_0/out vss 0.30577f
C1455 d0 vss 5.89103f
C1456 tmux_7therm_to_3bin_0/R1/m1_n100_n100# vss 0.10692f
C1457 tmux_7therm_to_3bin_0/buffer_8/in vss 1.28735f
C1458 tmux_7therm_to_3bin_0/buffer_7/in vss 0.74661f
C1459 tmux_7therm_to_3bin_0/tmux_2to1_3/XM5/G vss 0.55051f
C1460 tmux_7therm_to_3bin_0/R1/R1 vss 3.00001f
C1461 tmux_7therm_to_3bin_0/tmux_2to1_3/B vss 0.41874f
C1462 tmux_7therm_to_3bin_0/tmux_2to1_2/XM5/G vss 0.55051f
C1463 tmux_7therm_to_3bin_0/tmux_2to1_1/XM5/G vss 0.55051f
C1464 vin vss 23.7852f
C1465 comp_p_6/tail vss 1.09633f
C1466 comp_p_6/latch_right vss 3.49372f
C1467 comp_p_6/out_left vss 3.20258f
C1468 comp_p_6/latch_left vss 3.68918f
C1469 comp_p_5/tail vss 1.09613f
C1470 comp_p_5/latch_right vss 12.23842f
C1471 comp_p_5/out_left vss 2.08667f
C1472 comp_p_5/latch_left vss 10.47837f
C1473 comp_p_4/tail vss 1.56897f
C1474 comp_p_4/latch_right vss 5.50989f
C1475 comp_p_4/out_left vss 5.17613f
C1476 comp_p_4/latch_left vss 6.03696f
C1477 comp_p_3/tail vss 1.09611f
C1478 comp_p_3/latch_right vss 3.5009f
C1479 comp_p_3/out_left vss 2.06137f
C1480 comp_p_3/latch_left vss 10.47733f
C1481 comp_p_2/tail vss 1.56898f
C1482 comp_p_2/latch_right vss 5.48656f
C1483 comp_p_2/out_left vss 5.16723f
C1484 comp_p_2/latch_left vss 11.49738f
C1485 comp_p_0/tail vss 1.56897f
C1486 comp_p_0/latch_right vss 12.84132f
C1487 comp_p_0/out_left vss 5.23391f
C1488 comp_p_0/latch_left vss 6.03535f
C1489 comp_p_1/tail vss 1.09611f
C1490 comp_p_1/latch_right vss 3.49227f
C1491 comp_p_1/out_left vss 2.0627f
C1492 comp_p_1/latch_left vss 10.47733f
C1493 comp_p_0/vinn vss 6.06348f
C1494 comp_p_2/vinn vss 4.46291f
C1495 comp_p_3/vinn vss 7.44892f
C1496 comp_p_4/vinn vss 4.49649f
C1497 comp_p_5/vinn vss 7.17599f
C1498 comp_p_6/vinn vss 8.16656f
C1499 comp_p_1/vinn vss 8.11402f
C1500 vref vss 4.25902f
C1501 vbias_generation_0/bias_n vss 2.63421f
C1502 vbias_generation_0/XR_bias_4/R1 vss 1.61917f
C1503 vbias_generation_0/XR_bias_3/R2 vss 1.9113f
C1504 vbias_generation_0/XR_bias_2/R2 vss 1.5274f
C1505 comp_p_6/vbias_p vss 22.48268f
.ends

