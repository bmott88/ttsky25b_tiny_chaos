* NGSPICE file created from res_ladder_vref_lvs.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_6G5R54 B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_1p41 l=1.41
.ends

.subckt res_ladder_vref_lvs ref0 ref1 ref2 ref3 ref4 ref5 ref6 vref vss
XXR1 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR2 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR3 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR12 vss ref6 vref sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR4 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR5 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR6 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR7 vss ref0 vss sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR8 vss ref0 vss sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR9 vss ref6 vref sky130_fd_pr__res_xhigh_po_1p41_6G5R54
.ends

