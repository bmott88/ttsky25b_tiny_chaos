* NGSPICE file created from inv_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_PJMNR4 D S G VSUBS
X0 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 D S 0.16211f
C1 G S 0.02545f
C2 G D 0.02545f
C3 S VSUBS 0.11273f
C4 D VSUBS 0.11273f
C5 G VSUBS 0.31312f
.ends

.subckt sky130_fd_pr__pfet_01v8_MTNEXU D S G w_n109_n300# VSUBS
X0 S G D w_n109_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 G S 0.02934f
C1 G D 0.02934f
C2 S D 0.32105f
C3 G w_n109_n300# 0.1061f
C4 S w_n109_n300# 0.01071f
C5 D w_n109_n300# 0.01071f
C6 S VSUBS 0.18669f
C7 D VSUBS 0.18669f
C8 G VSUBS 0.22337f
C9 w_n109_n300# VSUBS 0.3924f
.ends

.subckt inv_extracted vdd vout
XMn vdd vout vdd VSUBS sky130_fd_pr__nfet_01v8_PJMNR4
XMp vdd vout vdd Mp/w_n109_n300# VSUBS sky130_fd_pr__pfet_01v8_MTNEXU
X0 vout vdd.t2 vdd.t3 VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X1 vout vdd.t0 vdd.t1 Mp/w_n109_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=0 l=0
R0 vdd.t0 vdd.n3 556.59
R1 vdd vdd.t0 547.24
R2 vdd.t2 vdd.n2 381.413
R3 vdd vdd.t2 372.113
R4 vdd vdd.t1 111.784
R5 vdd vdd.t3 79.0672
R6 vdd.n3 vdd 9.35164
R7 vdd.n4 vdd 9.3005
R8 vdd.n1 vdd 5.0275
R9 vdd.n5 vdd 2.53885
R10 vdd.n2 vdd 0.387074
R11 vdd.n4 vdd 0.381385
R12 vdd.n3 vdd 0.203152
R13 vdd.n0 vdd 0.106981
R14 vdd.n6 vdd 0.102352
R15 vdd.n2 vdd.n1 0.0996379
R16 vdd.n0 vdd 0.0996379
R17 vdd.n5 vdd.n4 0.0979576
R18 vdd vdd.n6 0.0937203
R19 vdd.n1 vdd.n0 0.0414483
R20 vdd.n6 vdd.n5 0.0407542
R21 vout vout 5.09101
R22 vout vout 2.59568
C0 vdd Mp/w_n109_n300# 0.01822f
C1 vout vdd 0.17246f
C2 vout Mp/w_n109_n300# 0.01232f
C3 vout VSUBS 0.36321f
C4 vdd VSUBS 0.88642f
C5 Mp/w_n109_n300# VSUBS 0.3924f
.ends

