* NGSPICE file created from inv_lvs.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_PJMNR4 D S G VSUBS
X0 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_MTNEXU D S G
X0 S G D w_n109_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt inv_lvs vdd vout
XMn vdd vout vdd VSUBS sky130_fd_pr__nfet_01v8_PJMNR4
XMp vdd vout vdd sky130_fd_pr__pfet_01v8_MTNEXU
.ends

