* NGSPICE file created from res_ladder_vref_extracted.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_6G5R54 B R1 R2
X0 R1 R2 B sky130_fd_pr__res_xhigh_po_1p41 l=1.41
C0 R2 R1 0.06364f
C1 R2 B 0.77617f
C2 R1 B 0.77617f
.ends

.subckt res_ladder_vref_extracted ref0 ref1 ref2 ref3 ref4 ref5 ref6 vref vss
XXR1 vss ref6 ref5 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR2 vss ref4 ref5 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR3 vss ref4 ref3 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR12 vss ref6 vref sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR4 vss ref2 ref3 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR5 vss ref2 ref1 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR6 vss ref0 ref1 sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR7 vss ref0 vss sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR8 vss ref0 vss sky130_fd_pr__res_xhigh_po_1p41_6G5R54
XXR9 vss ref6 vref sky130_fd_pr__res_xhigh_po_1p41_6G5R54
R0 ref6.n0 ref6 8.64891
R1 ref6.n1 ref6 8.64891
R2 ref6.n2 ref6 8.64891
R3 ref6.n2 ref6.n1 0.147491
R4 ref6.n1 ref6.n0 0.147491
R5 ref6 ref6.n2 0.0412986
R6 ref6.n0 ref6 0.0412986
R7 ref5.n1 ref5 8.6036
R8 ref5.n0 ref5 8.6036
R9 ref5.n1 ref5.n0 0.147491
R10 ref5 ref5.n1 0.0412986
R11 ref5.n0 ref5 0.0412986
R12 vss.n107 vss.n1 5255.26
R13 vss.n45 vss.n40 5255.26
R14 vss.n103 vss.n102 3882.06
R15 vss.n102 vss.n3 3882.06
R16 vss.n96 vss.n8 3882.06
R17 vss.n96 vss.n9 3882.06
R18 vss.n88 vss.n87 3882.06
R19 vss.n88 vss.n12 3882.06
R20 vss.n82 vss.n14 3882.06
R21 vss.n83 vss.n82 3882.06
R22 vss.n77 vss.n20 3882.06
R23 vss.n77 vss.n21 3882.06
R24 vss.n67 vss.n24 3882.06
R25 vss.n67 vss.n66 3882.06
R26 vss.n62 vss.n61 3882.06
R27 vss.n61 vss.n27 3882.06
R28 vss.n55 vss.n34 3882.06
R29 vss.n55 vss.n32 3882.06
R30 vss.n49 vss.n48 3882.06
R31 vss.n48 vss.n37 3882.06
R32 vss.n107 vss.n3 1373.21
R33 vss.n8 vss.n5 1373.21
R34 vss.n103 vss.n5 1373.21
R35 vss.n104 vss.n103 1373.21
R36 vss.n91 vss.n12 1373.21
R37 vss.n91 vss.n9 1373.21
R38 vss.n93 vss.n9 1373.21
R39 vss.n93 vss.n3 1373.21
R40 vss.n86 vss.n14 1373.21
R41 vss.n87 vss.n86 1373.21
R42 vss.n87 vss.n11 1373.21
R43 vss.n11 vss.n8 1373.21
R44 vss.n21 vss.n17 1373.21
R45 vss.n83 vss.n17 1373.21
R46 vss.n84 vss.n83 1373.21
R47 vss.n84 vss.n12 1373.21
R48 vss.n71 vss.n24 1373.21
R49 vss.n71 vss.n20 1373.21
R50 vss.n74 vss.n20 1373.21
R51 vss.n74 vss.n14 1373.21
R52 vss.n65 vss.n27 1373.21
R53 vss.n66 vss.n65 1373.21
R54 vss.n66 vss.n23 1373.21
R55 vss.n23 vss.n21 1373.21
R56 vss.n34 vss.n29 1373.21
R57 vss.n62 vss.n29 1373.21
R58 vss.n63 vss.n62 1373.21
R59 vss.n63 vss.n24 1373.21
R60 vss.n43 vss.n37 1373.21
R61 vss.n43 vss.n32 1373.21
R62 vss.n58 vss.n32 1373.21
R63 vss.n58 vss.n27 1373.21
R64 vss.n49 vss.n36 1373.21
R65 vss.n50 vss.n49 1373.21
R66 vss.n50 vss.n34 1373.21
R67 vss.n45 vss.n37 1373.21
R68 vss.n47 vss.n46 772.891
R69 vss.n47 vss.n33 772.891
R70 vss.n56 vss.n33 772.891
R71 vss.n57 vss.n56 772.891
R72 vss.n57 vss.n28 772.891
R73 vss.n64 vss.n28 772.891
R74 vss.n64 vss.n22 772.891
R75 vss.n72 vss.n22 772.891
R76 vss.n76 vss.n72 772.891
R77 vss.n76 vss.n75 772.891
R78 vss.n75 vss.n16 772.891
R79 vss.n85 vss.n16 772.891
R80 vss.n85 vss.n10 772.891
R81 vss.n92 vss.n10 772.891
R82 vss.n95 vss.n92 772.891
R83 vss.n95 vss.n94 772.891
R84 vss.n94 vss.n4 772.891
R85 vss.n106 vss.n4 772.891
R86 vss.n105 vss.n1 686.553
R87 vss.n40 vss.n39 686.553
R88 vss vss.n42 341.459
R89 vss.n42 vss.n41 341.459
R90 vss.n108 vss.n0 341.459
R91 vss.n108 vss 341.459
R92 vss.n38 vss.n35 252.236
R93 vss.n44 vss.n38 252.236
R94 vss.n54 vss.n53 252.236
R95 vss.n54 vss.n31 252.236
R96 vss.n60 vss.n30 252.236
R97 vss.n60 vss.n59 252.236
R98 vss.n69 vss.n68 252.236
R99 vss.n68 vss.n26 252.236
R100 vss.n78 vss.n19 252.236
R101 vss.n79 vss.n78 252.236
R102 vss.n81 vss.n18 252.236
R103 vss.n81 vss.n80 252.236
R104 vss.n89 vss.n13 252.236
R105 vss.n90 vss.n89 252.236
R106 vss.n98 vss.n97 252.236
R107 vss.n97 vss.n7 252.236
R108 vss.n101 vss.n100 252.236
R109 vss.n101 vss.n2 252.236
R110 vss.n45 vss 117.001
R111 vss.n46 vss.n45 117.001
R112 vss.n41 vss.n36 117.001
R113 vss.n51 vss.n50 117.001
R114 vss.n50 vss.n33 117.001
R115 vss vss.n43 117.001
R116 vss.n43 vss.n33 117.001
R117 vss vss.n58 117.001
R118 vss.n58 vss.n57 117.001
R119 vss.n52 vss.n29 117.001
R120 vss.n57 vss.n29 117.001
R121 vss.n63 vss.n25 117.001
R122 vss.n64 vss.n63 117.001
R123 vss.n65 vss 117.001
R124 vss.n65 vss.n64 117.001
R125 vss.n23 vss 117.001
R126 vss.n72 vss.n23 117.001
R127 vss.n71 vss.n70 117.001
R128 vss.n72 vss.n71 117.001
R129 vss.n74 vss.n73 117.001
R130 vss.n75 vss.n74 117.001
R131 vss vss.n17 117.001
R132 vss.n75 vss.n17 117.001
R133 vss.n84 vss 117.001
R134 vss.n85 vss.n84 117.001
R135 vss.n86 vss.n15 117.001
R136 vss.n86 vss.n85 117.001
R137 vss.n11 vss.n6 117.001
R138 vss.n92 vss.n11 117.001
R139 vss.n91 vss 117.001
R140 vss.n92 vss.n91 117.001
R141 vss.n93 vss 117.001
R142 vss.n94 vss.n93 117.001
R143 vss.n99 vss.n5 117.001
R144 vss.n94 vss.n5 117.001
R145 vss.n104 vss.n0 117.001
R146 vss vss.n107 117.001
R147 vss.n107 vss.n106 117.001
R148 vss.n105 vss.n104 99.5008
R149 vss.n39 vss.n36 99.5008
R150 vss vss.n44 89.224
R151 vss.n41 vss.n35 89.224
R152 vss.n51 vss.n35 89.224
R153 vss.n53 vss.n51 89.224
R154 vss.n44 vss 89.224
R155 vss vss.n31 89.224
R156 vss vss.n31 89.224
R157 vss.n59 vss 89.224
R158 vss.n53 vss.n52 89.224
R159 vss.n52 vss.n30 89.224
R160 vss.n30 vss.n25 89.224
R161 vss.n69 vss.n25 89.224
R162 vss.n59 vss 89.224
R163 vss vss.n26 89.224
R164 vss.n26 vss 89.224
R165 vss.n79 vss 89.224
R166 vss.n70 vss.n69 89.224
R167 vss.n70 vss.n19 89.224
R168 vss.n73 vss.n19 89.224
R169 vss.n73 vss.n18 89.224
R170 vss vss.n79 89.224
R171 vss.n80 vss 89.224
R172 vss.n80 vss 89.224
R173 vss.n90 vss 89.224
R174 vss.n18 vss.n15 89.224
R175 vss.n15 vss.n13 89.224
R176 vss.n13 vss.n6 89.224
R177 vss.n98 vss.n6 89.224
R178 vss vss.n90 89.224
R179 vss vss.n7 89.224
R180 vss vss.n7 89.224
R181 vss vss.n2 89.224
R182 vss.n99 vss.n98 89.224
R183 vss.n100 vss.n99 89.224
R184 vss.n100 vss.n0 89.224
R185 vss vss.n2 89.224
R186 vss.n42 vss.n40 34.4123
R187 vss.n48 vss.n38 34.4123
R188 vss.n48 vss.n47 34.4123
R189 vss.n55 vss.n54 34.4123
R190 vss.n56 vss.n55 34.4123
R191 vss.n61 vss.n60 34.4123
R192 vss.n61 vss.n28 34.4123
R193 vss.n68 vss.n67 34.4123
R194 vss.n67 vss.n22 34.4123
R195 vss.n78 vss.n77 34.4123
R196 vss.n77 vss.n76 34.4123
R197 vss.n82 vss.n81 34.4123
R198 vss.n82 vss.n16 34.4123
R199 vss.n89 vss.n88 34.4123
R200 vss.n88 vss.n10 34.4123
R201 vss.n97 vss.n96 34.4123
R202 vss.n96 vss.n95 34.4123
R203 vss.n102 vss.n101 34.4123
R204 vss.n102 vss.n4 34.4123
R205 vss.n108 vss.n1 34.4123
R206 vss.n46 vss.n39 15.286
R207 vss.n106 vss.n105 15.286
R208 vss.n109 vss 8.75059
R209 vss.n109 vss 8.6036
R210 vss.n110 vss 0.831056
R211 vss vss.n110 0.774111
R212 vss vss.n108 0.489974
R213 vss.n110 vss 0.231056
R214 vss.n110 vss 0.174111
R215 vss vss.n109 0.0632894
R216 vss.n110 vss 0.0135208
R217 vss.n110 vss 0.0135208
R218 ref4.n0 ref4 8.64891
R219 ref4.n1 ref4 8.64891
R220 ref4.n1 ref4.n0 0.147491
R221 ref4 ref4.n1 0.0412986
R222 ref4.n0 ref4 0.0412986
R223 ref3.n1 ref3 8.6036
R224 ref3.n0 ref3 8.6036
R225 ref3.n1 ref3.n0 0.147491
R226 ref3 ref3.n1 0.0412986
R227 ref3.n0 ref3 0.0412986
R228 vref.n0 vref 8.75059
R229 vref.n0 vref 8.6036
R230 vref.n1 vref 0.831056
R231 vref vref.n1 0.774111
R232 vref.n1 vref 0.231056
R233 vref.n1 vref 0.174111
R234 vref vref.n0 0.0632894
R235 vref.n1 vref 0.0135208
R236 vref.n1 vref 0.0135208
R237 ref2.n0 ref2 8.64891
R238 ref2.n1 ref2 8.64891
R239 ref2.n1 ref2.n0 0.147491
R240 ref2 ref2.n1 0.0412986
R241 ref2.n0 ref2 0.0412986
R242 ref1.n1 ref1 8.6036
R243 ref1.n0 ref1 8.6036
R244 ref1.n1 ref1.n0 0.147491
R245 ref1 ref1.n1 0.0412986
R246 ref1.n0 ref1 0.0412986
R247 ref0.n0 ref0 8.64891
R248 ref0.n1 ref0 8.64891
R249 ref0.n2 ref0 8.64891
R250 ref0.n2 ref0.n1 0.147491
R251 ref0.n1 ref0.n0 0.147491
R252 ref0 ref0.n2 0.0412986
R253 ref0.n0 ref0 0.0412986
C0 ref5 vref 0.06887f
C1 ref4 ref2 0.06887f
C2 ref3 ref4 0.00359f
C3 ref6 ref4 0.06887f
C4 ref5 ref3 0.06887f
C5 ref6 ref5 0.00359f
C6 ref6 vref 0.19117f
C7 ref1 ref0 0.00359f
C8 ref1 ref2 0.00359f
C9 ref0 ref2 0.06887f
C10 ref1 ref3 0.06887f
C11 ref3 ref2 0.00359f
C12 ref5 ref4 0.00359f
C13 vref vss 2.14919f
C14 ref0 vss 2.42437f
C15 ref1 vss 1.54901f
C16 ref2 vss 1.48014f
C17 ref3 vss 1.48014f
C18 ref4 vss 1.48014f
C19 ref5 vss 1.48014f
C20 ref6 vss 2.23319f
.ends

