magic
tech sky130A
magscale 1 2
timestamp 1761320183
<< error_s >>
rect 384 843 442 849
rect 384 809 396 843
rect 384 803 442 809
rect 384 315 442 321
rect 384 281 396 315
rect 384 275 442 281
rect 384 196 442 202
rect 384 162 396 196
rect 384 156 442 162
rect 384 -114 442 -108
rect 384 -148 396 -114
rect 384 -154 442 -148
use sky130_fd_pr__nfet_01v8_PJMNR4  Mn
timestamp 1761320183
transform 1 0 413 0 1 24
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_MTNEXU  Mp
timestamp 1761320183
transform 1 0 413 0 1 562
box -109 -300 109 300
use sky130_fd_pr__nfet_01v8_MH3LLV  XMn
timestamp 0
transform 1 0 158 0 1 257
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_TMVPE9  XMp
timestamp 0
transform 1 0 527 0 1 213
box 0 0 1 1
<< end >>
