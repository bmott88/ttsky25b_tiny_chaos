magic
tech sky130A
timestamp 1761410844
<< end >>
